PK                      archive/data.pklFB ZZZZZZZZZZZZZZ�ccollections
OrderedDict
q )Rq(X
   fc1.weightqctorch._utils
_rebuild_tensor_v2
q((X   storageqctorch
FloatStorage
qX   0qX   cpuqM tqQK K@K�q	KK�q
�h )RqtqRqX   fc1.biasqh((hhX   1qhK@tqQK K@�qK�q�h )RqtqRqX
   fc2.weightqh((hhX   2qhM  tqQK K�K@�qK@K�q�h )RqtqRqX   fc2.biasqh((hhX   3qhK�tq QK K��q!K�q"�h )Rq#tq$Rq%X
   out.weightq&h((hhX   4q'hM tq(QK KK��q)K�K�q*�h )Rq+tq,Rq-X   out.biasq.h((hhX   5q/hKtq0QK K�q1K�q2�h )Rq3tq4Rq5u}q6X	   _metadataq7h )Rq8(X    q9}q:X   versionq;KsX   fc1q<}q=h;KsX   fc2q>}q?h;KsX   outq@}qAh;Ksusb.PK�od�p  p  PK                      archive/data/0FB ZZZZZZZZZZZZZZZZx�-= �<�q� o���=@/z�?S��K��=�������<���=��(���!���96��<:�.>7F��3?|ο� �?�=�?*-���]f?��?ծ¿��S��,��$E^?�"����#]�i��<F���Z0>&Z��_u��{G=�� ��>�w�I\?�{����=��4>�J��ٌ>�uȿ"��>?��њ�>�ئ��ف?{ϛ�Ww�>�.�>�J.?������������ž;��&��s�dE�>�W��y^�}�>�Z8�=�,K����<����z�u����Ѳ���.�Z�@> ����ᪿ������ž�����5�2 ��l2�~dz>�g�H-�=�����`��>6[�=�Ȓ�U%�F?�=Mk��#�g�D������?��;��x��_Dξ�'���B�3B��=&L2=����0���S*���{T�����܃�凾zM�>�u�����>C[��?���>����n�?#�.?��?��]�f��H?q6����?(?���?l��>�S^?�N�":�>C�P���u>A�?��X>�=e?.�?+���ws���#�0�B>^\���	��`����������H>Y<�a��;�)����	�:��>L[R��>𿆳a��||>_��;�?��ɾT 1��Q<?�t:?�����=�������ؤ�M����?�/>r�>��}=p=>�-�>K�L���M?�ą?"w?�<�>�i�8�/?��]?u�?lR#@<��?��O�\���l���h����
���'�D6��������Y>�Ɩ���>(���7>���<�����y�>[�ҽW*ɽ��/�m��Cy��<���O�>>)�<'Rg>�f{�:4^��R�'�L�o��=�q����?E��>�+%>r]"?`�+��&���'?���>���Ԛ}���Z����>8�=^,���'�?�k?�
*�N��=D]=���<{�9���d>e\l=�CÉ��!>�����þ���Zr�=��H> �>c�5?1��?��9?k��m�>?`�ξ��R?9���*�?:��Z�x�����w�?��?��W�e7 �~"������ۖT?���λP��8?1�w��SĿ�1i�&"�������Z�>�t?�~*?�p�(Ѫ��?�x'��%?��Y?$Ʃ>�鞾�:�<�C�>�����Am��Զ��(��)�E>��<�d&��%�?)`p���8W�Jf���m�<f��4"|����?��˿3b���K��.t?5`O��`"�%�P��w&�0\B>���=S�1=�
��j�>��<��H��W���e[z�ќ��ՙ&�/=$=�<@��(���j�/��'b��6<��<R?��?�2.=�r�?B�?��l?�;�>�@?�+?���?C�"?��6��Ψ�
f�=LCd��';?v�?�o�>�{>���5�k� ?���?��`���	�����@C�>5�⿶����^�F+J=g�r?�#@��xk�J�澽k�=9��]�a��3,�/9b�z��=�6}�FYŽ�	���>#�.�\��>�4������K���m�>
:�?,gR�Oi�cR�O�?W��3�����9>�?��ѿhOa�⾾l>��?�N?������l��ʾ�Rǿ1���l�*�a���:?=?��b=��R?�+*�;�پf-���aſ:�ž�g
�M������H�@��?\[�<�X�?�G�>�?cv$�5�>6�>��ai5>���?�U?�Vb?,C�g�&?58b<��t?\}��+P������$B��n�W�g�|c��?y_���2?r�z>�q+���ӿ��Z��;?nw��y��?tP����>�,޿��п]�>C��>t�N��5=�>㾿>`���:o�bpоȮ����K���<���ľlaR��"��o�<�L?��>�v`�������>�0��ю��ׁ�>P�G�Ļp>�h����O��=x��.�>D��>�꪿)X�[�=�R��{6�>���s��Z�T?ΰW�Q�9���_����>;��>V���>�⹾�mX�у��G��B܈?�Pb?���<���i=�~���c��Ü�mV>�,=��Կ�7���aʾcq;?Ī=[��?�{�$"�>#-?򠘾WG,?S�G?�=?uqZ?�g�Z���X>'��$��>x�?rۿ��<0G����A��Î�c$��wU��a^����K�[?��e>���Sը�¯ؾն��� ;?���>�?��> 9b?��ҿ��@:�?�r9>�(?��'?�? A?���?p�?)�?�?�bx�@O�>"Wh��u�l˞��M?��M~�����ۖ?(���Y�>efd�8H�=�PI�\V��S�z<>�0û��S>��G<F�f�J#u����@�Y=�a9��4����*����8� ���%��pG�2
>�+&<% a����)�j?�z>`:ſ��?���'W��@�|�a6�?��KB鿧_u?�����+�>j��=j����0F�ud�?�z�Ҩ?�mh?8�R?|&�?A2�?_��>I�6?'�4?� j<�@�5�?R;?��G?�>S�����m��r�?�m��.�ګ���T��g�
�$����\�H�W����Ԟ��̽pT�ă�=�vP=�� ���p��<��K= ��<@��k}���]��Z>����`��=���v笿f���:�?�,��Ԇ����f�uLƽ����n?�k���D�ю!��lV�滛��!��$e��m��?�@�> 3? O>+�?O���Y�C�= ?Ȅ�u�r��9?�_#@���?�".@1m?|�?�(!�kT��]*0�6ǿ|r��� �j"�|t!����b?V�>��~�{ ���@�2����A�]v�:�Y��94>���=	ᇾT�F���~���~�*��!kW>#X�7�<�C�=��*�O�=��r�s �:�5�!�6�=���u��v��R�>	����d=V�=!-��jV$��? ž�i���ֿjO���C=N�m>���W?��b?��?Ka7?Ä�}�����?�㌾��3�=���U��n�>��=-�:��\�>��[??,@�d�տ�cN�?�нcw���k7�>��-?��ĿMM���刾�P�?�f*?ژ�>ƹ>�#��n ?I��?:�>�{�s1�>p���AW����=�1�>�E>�<���6��־�<?�l��T�C���>��b?J�ؿ)7Կ���M>?n��>��ʾ>������3ݫ�h�(���վ<rO?�����3�/����� ��� @ͿȾ�c�>u�ǿ<�?P�����	|2? Z>4�T��[�k$&�Pq��ݾXX�������R?��>/�u?���=��[>��ݾ� �>���?`�����=������^?�Ͽ	ʡ>_M�=�����Lý���>�kb?�G�B�Y?��� ���i����@@� �a��yG���!7?8	�Lt �b*D?(p/>����4t�?\�O�5�(�į���.�"�2��]�?�2�=�ҥ�Zga�p����S=3��=&��=��9> 7��e�=��I�֖'>aZ��Y�ܲ������ �н�k�@DD�����m�?D��� ����? ���'��3�e���ྦ�67�=�ǋ�����=,�?�A�7�>1S�>9��M:?�<�6td�r�>YW�>�R�&�:>�??+����f�/��ҴM?��>��~>�=�LD�	?���<3�J?u�?��?��>�O �c�?f^P�����ۿ�������p>���TԻ��Z���7��3��+w)?��C��S?#��g ���d�<�Q����+4�1���mhž�wɾ�W9�MW?��>%�Q>4��>�G
��R��e�>Ymh�r�0��B龘�qm�x�J���ʕ����>��#���ξ���>��+�L��>lQ���;z>ƅ;��q��ޚ�=���>E~?�a��N���̮�GK�?���>)*������H�>!�C�&��u.�>6s�>���:���w?�4��ӹg?g��?� �=�����7��9Q?��K?U��;~� C?����q���H���?PK7�C�      PK                      archive/data/1FB  O�K�NR�'��3�;�l�'���?|c��Tq���'�߽���u_>Ӣ�(�Z�B3N?�������=����b?��?�O0��,C�+�>�%9����>��Z�����_�=��@��/����ž�����'?f��>  >�ྒw�������>f��Q-6�*.=�i~��;�c"�=s"� Ͽ��T?==}>��>>]���U=�I?3e��B�>zԊ�	�,�p�V?7+���NE����?g����0?�ń�PKp��b      PK                      archive/data/2FB  |5�=�>=�vE�o�=��<����ȼ�i_=�����t=�{��?������?���Z�C��=Q9�J�@=l�彦���&4��/��J�=@4���e��S;� ��q"U��]l���=E���+����������$�w�� t�*���ܜ�9/+�`hܻ��=�͆=�˵<褃�;0���$��װ���D=�'$�?x��s�&t�<��E�v3=x/�������"�T��<[�<s,�\Q��A�f��=a�I�V� \�������M���̽
u���Q=2����<��<; ���{�����<��k�V�%A���=��=�Z=h�i��*��"Ҽ�@=Jo�=E�c��_����=��/�r�ý���Ƀ��+=�R�U���ؽ�V�����i���g <v󔽶4ɽ@���GP��ꊓ��
�������*# �_��(g7�������<����t�= D��؀���<�
O=t=ĽA���_7��Ľ����-������ǻW#����/&���g=C���U �������^z����=b�L=��=�{|=�EW����r����=�zd;N���`7��F�p��Y����<��|=�_�<v���F=h�$�"���#���f!�ۈG;`T�</<Kw=�����虼e]���̑i�h;�������ϻW����|�<�A��iǽG6K<u���h$d=��`<�z��cW!=�ϼ�uѼ�W��,I��.�q=�@�� .��L��0?�~��>x=?�-�?PV��N�>�x������+����>�A?<�����B�*a�X�>r@�ӈX>��=��	ux�p7h��>�����>Z�o����O*��#�?9[�?�q�%
�=��(Yս��ֿ=��D�+=�$��ɏ����@���<��"����8���l�N���؏?�
����������X�J#�>���=+�i�>2����?~A��n���P�?�딿V�+?�6X�2j�=K�;>�ܜ>�ǿu�O��a�-��?A.9?u����f�f�_����g2������9?��!?����ջ�<֪*>��a� >T�����@����=ʽ!��?D�w?'�����)��ွ��=?,?Uצ>�U�<����@���(�'�|"T�Fi��M����?P_��*��>5(�_?��7��@@�mݾ�ľ�j��M���6>Pz'�L@�=��Ľ�`��#�����Wu�Ů�>~6����>v����$�c=���=��<J��9�O�@j�=���<��M��׻�T=�&��W�=�.��Y+��Cӽ4:m�#���Pؽ��꽨�o�X�<���7r ����|���|gr=��+=}O�U�< �|��O=rA/���8�|๽�KZ=�E����ֽ1Z�`��=Rk � ��<plu=�`S=D�����=��ܽ��7�;���8�<�7�<}��ԟ=!̮<̀/���=jT'�)|����O=6+�4)ļ4f�<�F���ƽ�1�=*�S>��>��N�ߣ�e$վ�����?�Ϳ��>��?D����?Yu���I���N<���^�m?��� ��ā>�����?c�ο�0?R�$?�6��0f����'?��L?� �>��ֿ@�>Ho�̫_�l;>Լ�?�2<>腍��[?�7;=H9�fd�6�{��<��n�h 5��Ŀ��m?>��>�e���ľ�m=W]�?겨;��=b���*?��j>ߝ������Ҿ�,��L�h��#��`��>8��6�=��Z�=ȱ>u�]�!��1�>���S�F�>F+E>�9=Wp�<��3�F?�S�����m=�}�\0��y<��k>p��!'�=�����ῳ� ����<0�P>}`f��G�>.�̽40Ǿ{�0��ѽ�r��ܣ�<��"��#�=e�y�!!Կ*ν=E��i���!>�Z��">��⾿�ľ�o>E�R�b���2����k���G����=�o^�|�翢����=F�ῌ��~����M"?T8���N��އ>k5��{�>=�>)z_�M�P=���>P�<�f�>{"о�೾��.>��F���<���?x,��c�=^,?0��>�#��!X������Y�uj���:$����Yl? ��9�5��Ŀ�=�þI����#�d��=��?�)���?������Qk&�w�
>E�f>6���T&���a>�\	?�8[�|�D=���?���;���x/��?Hi>?Z\�=6�?&亽��]?Xg�?6��?IY��6�F?R���V矼y��>�u?���i�>�<4?�lj�#�)���%��J_��!��1�<��Z>�G�����?N�>���Y�W���y�K�N?��=��?H�#>������C��>(?�=x\����p9>>����󢿋TK�˛=�q�*����4A?�����)�&�W�}2������1� Y?�)��0c)����=��?�: ����>s��?��
��L>��/��0��^���Xe�=d�?�o�>1BV?/e���xQ?$����^�>��?�C�t��>�m?�奾��> @��?P'��=U�=lyh�eX�>��c?K�b��|>|_w<��?�֮��QY?U�?? %�?#�>g�>":;\�������˼d䒿�ך�`]@V�I�꾀D��$S�?�>�=���/I�>�#ʿ��N�:@�A?�Lg?�>4?�5�?���������?3���Jv?��-?�����b���b����=Il��G:?���^k����˽�#�����?y6��T�U����¾�+����>!�>�N��o/?L�>�)?�/=ޓA��+ؿ@ͻ?a?�A�?���=W����,��3H�?�.�>L��>��?���>G�i?;�|��Ms??�8��=�C?J(#�_c�^�ٽg�8>i:v�ދG�`���u �(J�����p����.@��>�j:?��݌	�4�5�I���Uc<�"��&�}? ,����>�-u�]���/&b<���Y�>��;�d��q�)=2h�>��M=�C�u������=2��~���.������*k�=�޿Mq�>���k�D���L=t��b����5�=����N�S!k=�����>���?n%�&�ݾ�0V>��1����̥�x��<�]>��W>Y���͞=��4f����N��ݣ=}&�;Z؄���Ѽ�d���5l�1�>bq����=x�켴T�=Nqe��-�1>�	���Aބ��վ}K#���5V̿=�l?d��=�+	?�)��q�I>ӱf?�
��C�>*�j?Q��{>�5?*��2�>W��P��~'���ǿ���=<��x�O�36��s=�V�?��������P�>q�7?Ҵ=e$�?�	=�k	>���1�>��B>qX�����\"?&,����_�?Ȏ=[���嬿z����8�!�?�����$��^G?e�?���̂�Q����O�%62>N�?Tw7�@?a�Z?��޼�|	=�%�=eI��D'X=ft�<�)=3�5�\�>������v�}����U&=|<� ��3ܼ�*����p�� �ҽh�k���<�G|=�|��g1�E��M�ʽB����g=��"�������b=t��R<�>�߽��I�,���|����"�z5�=��=h��<�,I=�$W<��q���=Y�۽Pͽ����j=�)�����l=��������b��<���;���;f崽Y"�<-"+�/�Ž1N���	�;k����|?���>�A�=V�C�_��X�?o��m�>�l
?2_3��,�>�0�>E<P��6=fR��$F?24�EN���8>·�s����(��hF?��>�kG>d�ݿ��3��>�>�ǉ?vD?u����x?j�%?��A���>=%�?�����O�>�[�<4�k�����y?/J��E��2�7>܂���n��"xQ�%W�?}(ƿ{-�L̵?���x��=e��>��ͤH�ʞ�>�V6>H�¾�-*?櫳��>�G�>��S��\>��J�_?�=*a�����z>�?����{h�>��>�{O�&�c>B�Կ���=���>��2�g�~>���J�|�D�>��~?������?�X%?���*^��?����G������MG�5B���'�
*;=�I��6�e���t�R�Lȿ���7��0@ <;2\�;�ӿ�w>x8@?�k� ���z?�>�띿�l|=��%�M?3�A��0}�S�=�1���S#��<���⽎B� �R�V>�U�=���f�x=�,Ž�Ҽ��{�%ռ9��Q�:$�=�Q���<����=:�=8�U<��=Ƽ��<�����3�J9�=y�½z.e�X9+=x3)�P���L޺�]�½�e�R����2��2νT�p=u����Kq<�佘�1�J�4�V��=t�/=�F����� �ɼ�U޽�>=��3�]ɑ�X��?��0 �=�k˽�Z���(�=�z����ƻt�e�����g=�چ�F� �=?�W�k�L?4	���̾1�2�A百�R�>l��=����H>ـD?���b�>+y�
�<���)>��;2��=YC��|�������!�#��>uJ�t����:I�!=�>��$�9���������8����v+~���=o��>A�b>L,��8A���|��V`�3�I>�j���f3�����ѽ���>@S<��:;�
kU��X��"ҽh���!��_���
�H��=�d��ѵ�+|�<0{(>>��L$��Op+?��H>�}n�Vg���!^�ޥ=?�|����>�G=Q�տ���>A�y>9]�-��>�?�~?~��\D(�L7>�B�ӗ�۶`>�����<�Y�W�Z�ܾ�򾐄�?dC>R�Ծv1������GaN���>گ���
L�$v"����+�O�Dg���v�d��=� A��bƿ�]?�ՎP?���?7 οl�8�U�ƿr��c#�=��̿ ��N���]P����E��>�z����>�׽�q�;�t��i�?�=h>�<��q?UQ�)^��(:>+cпդؼ���>�*>��i��q����V�-S�;�%�|����=���KZ���>>B�?g�=��̍K>tc�0F���̾ad�?h�m�Q�\?���=�P��h�>��M�g7J����>������=�?���c�uk:�J�=
 W?���}i/�[����i���?��LB�<{2þ�9���o/�����ĕ�]�{?�*���L?���h뿠	����A<r��=
Q��@o.�]��>�&��x�;<�%�=�ZI=�Qk=]�=bD#��N������:^=���<��5�.J}���=
�<�{a���d�����ܹ�z�½P��m��ZF�ص�O�v<�����|<J��UX��ն���Ki<��� o`��N��V=�$����������B=o���* "���~=&�7�	���:��5:<*�Ǽ@���}���ȼ�H����7L=M��=2ʽ;�$6�n�=� ���S�?�P�>|7?�x%>�y����靝��k�>#��H
��B�>g%?��q?#�>�<�ne�Q>>x��P%>�?ޔ�h��?�i�>��G�=��>�QE�p��6)�>J�>?�<¾g�>���>���1-�?n� �u5'<Tھh��>��w���I?���&?�e&�O5"�:=ȋ�`��������Yq�m�!?c��>ӄ�>mr|=h-,@���"�;��It?�(=�p? v��f���0V.=�O�;F =��C<��sn��k����.H�TԌ�!�=��=j�����<˗�<y��QAI<0nݽfjl�����Bʃ=e�ؽ�#=e��u[��$>�:lǽul<�!K�Gro��<s�2��^p�s�ɽ����l཭�����������G����<��=Z� ���/���8�
t�=5��A��9fL���L��s�<��A���ɽ�B��[��"�����ʽ~0>�n�B���ں�mk�T4�q�<9�� �<��Ͻ+�Y��}�nW����ǫ�=�:�}*�7�=c�<y�9ǒ��|ꮼ��J=�|νP�L��Ž~~��'>�`�<�6=��`<ü��(��Ľ���<k؄��R'�.b�=�㦼qF6=�o`�. �=~��9��W� �{<�1�<)�ϼR =\^>�X��$VV���;��=�5��¼ Av=s�n;颇�(����,���f%���<��=Hԧ=S��Ha����>s���x=�X�<�o��O�<X�����ֽ?���M�����4����RǼrV=xV���#"���=x'�� -��}�|���=@�н�%\:"~<j��;~Ԧ������X˽���偽�����;����/�=�w�<�̽�l�=t���� u��K��N�����s=�1��h"�g׻�6� �/:�ɯ���(���.<@�<�.�;�D�a� ߼m�
��F��b������E�u��-`<xɮ��lb���d��R�r��;�}=��c����А��?�_?.���ͱ�����?A�>�Z�?Ҽ?�׾��K*��O���~��s�>�n�>q���fiŽ��=?��>f���|�����V�?� �>C�)?�Pu�+ݾ���?�A�?5�>�H@�8��CU9����t�?=t1>�8�����>K�C��8�>"%�=�F�>��߾�����ؽ��z�<��3HZ�9X>7-*�����Agz>�m�?�<;�l�1��4U�$���r����?��E�X��>Lkн�U���\�����V?�ڟ���2?b*r�C	6?���#M�!��>��=�߿Ah	>�<?���E?�Q?JӾ?~?�j�<]��~+�9�i��>�@��z�?"׿�bȼ�@p��1�=�d��A#��Vpɽ�9U���=�mG�yi��[�=1�����!X:���g=7����>� u>x���~h��h�;�Կ�>��	�r�Q?B$�q҄�6kQ=�co>P��=��?��¿ʬ��t�Խ|� =Ӵ��XF�m��=<�D��@� ����>�51>������>+���B�>˄�?�Q鼶&�>|c?�rm���&>%/�����?���|���/>C��3���c�?�I?��.??���c������U�?��8?�v@�I��\Q>p�ؿ�2⾺>��F�=(а?yU����7?��O=������>V�l?��=�p9�=��>��G�)��,�?�a�?[?���|q@��2��	!�?*��ʿcg�?�+����0�i�F�)|&����<M�>�>sD!�:f��9�_׾Ɔ�W=��Ă<Ք��f��~���H>��ɿ˂>	�R����>W����=�z���"���5�0�?{=?����`!>�WR��⥾�?jѲ=�J?󃉿�_�>��)��D	���#?��==5�->��>�h�XP%�i��?�Qӿ/@`p��ĥ=��?󤖽�V�?��h�w�? ��>�K+>�Ƚ0�_<R�ﾥ�>���'��xJ���r����<��<��ֻm�<�>W0ռ���'S����N�,�)�˙B��*ҽ֯6�*Wѽ�&��X�����<c�»żI�!5{=�ǽv�<�Z#�U���o��޽��*=���U�
�t�ni�=b"��x��R�<��=
��<b<˽�ν�뽅��<����t=;E���;��ؼ����9�ٹ�� ��'wἾt���	��W�	���-��$��R�==�*=�3�.︔�ƽ�p`��=�����`1=�ʽ�ٽ�4��uw=�u=wu���"�Ň�����;���=���=������ؽYK�=G�D=��ݽ��ν�0�OT�ǤG=��ѽ���X�=�Ζ=�V��?���џ��.&�_[Q=� =�+�=d��ҖŽH��<��=FW��t=
n���9N=����z[=�/^<���r3ƽ�W�= �}:����8U��P�1���<�o�=�Q0�|Q������ȽV;��{˿=�!=��=�+��O����=m�e��؏�� �=E+8�X�;҇��yG>fy?:޾\�S='6�>b�꽁��=Ŗ"�]�9To�}���̍==�*���.?V�X>X �?�]齴n��	���u?N����p����/ʿ;�U���^��3$����A?̿ܿ�h�4���Na?O~���;դ<�ɜ?9p��67=�C�?�g�a`�����=�K*�g>ɩ?�lm��H.>t�ο/`>~��]�ٿF����>+�ֽVl����=|�I>2b�>M(�F�H��(�<t����=�9���J=�߉�yɼ=�}��k�'��y��)�<���=��̽�6c��p�;��=��vG��)���@�j��0L�{��=��@�t{q�*�G�g�����m=���$ ٽdA����1�l�!��� ���3<{K��b4i�(��1Ef��ܘ�W���W�=~�ｭo�h(p� �G���=�P��N����㎼� �Լ��Լ$����˽p�,=#^�k&�4�<
���7e<��={��0��<��=P�>B劾�9����<W�<���0?!��u!��#�AD;�m�� T��G�=@�\�S	��V	����$� �F��۽�F2��~�>�C��@�u��n?�^V��u�>=���=t�;�8s�o]�����<_e���>z�=�̽���>�0�N���G�|��b���#�0�=
�޽V��˩ɽ�2)�Y��=m*�?�֠=4I��N]��]5<�"��{پ�8�>U¿>�C��ӹ=�A���b��죽��e��[����I�������0�ݽ`���6��<��Ͻ��������A��ȼ��}����=�����;!��fe=]j��_=���d3��*�����g�����<�������׭�F\�<;�x�iF =�������0=���<Z�����2�pb�=�_��[3�U|i<�8�����)�g��=�		�}�=�܆��y=�^X<u��f��}�=f�<��<��<�&���KƼ�db�}���H+o=�����4?���Mf�m��O�>��
�Aj��.�>�gH?��i�>��;>��=4&3�ɾ`��ֽ���Ӿ��[?6{r>����;ȿv�>r�>I�d?�c??�$�W ֿ��l?�w?��:���	�?��3����o�h��7����B��@ ��r��d�=���K���HF=?��߽�`�a�ѿ��(�u�m����>�D7�e�=*@?F�2��Io�e4���%�� <��c?�mi����=@�6?]\�j����p������J���8?� ˾}p%�#ſד־y�>t)x>G'����>|��>T���f�>��->6Y�<�k�>��wJ>�z��[�?��cʽd/��J{>�n�>G�=bտ�y-?�I>e{�����׾�i>�R����ݿG�	=�����L�{|����=!🿩?r�KO/��4�=������ھ�����ؿחK>�"\���M>��޾u�"?�%�:y��?'P���5�/ۑ?�=�>�ܿ9���c�=ܣ=�Ӏ���q<D/>��=�/v��=/?��~�|��P����R�?�꨾��k=s��=�$�1�=0��>�_�>��οL��LY��6����ȿ��8?e?�#����=Aܿv��W��>xAX��@?<{�>ԓ�>��$�dz��h�p=�
�>���Tҿ�ք=[���U�Ծ0�0?���<��;��Կ�m����>�߽������?D=d��<�X[�<���?�/���<��o�?ˀ����L?��A�N`)������[$�g��?��
?�i�Ȅ�>�g?��:���
����>j|��@!�X�>���>b��E�u���Ŀr��=Sڿ��%��-z>������8���t5�2�/��8�?P�
��	b���+��Nh?,����==�^?�;*>���A�z�5�i+
��&��� ��`�:��o.?��~�O�I��Ĳ<:4����習���-?���ѿ�y4�,9�>����2;����Q=�H��	����z��q�>��E��Fz��M���n�>`��=A�(�{2=�8�=�����'�i����B�+埽^�=)��S���-:�=�r=������=9�ǽ�
��#��
�(=2=D=�[��x���R��u��R��T׼�텼�w��m�F<o��ʆ�Zl��3-�f��=˳;�GM��'�7=�D�	��p<ܼ�4�=�S���3F<�=$�!=�`޽���=�e��>Խ+N�=\�ѽ]��/���4��=�|���ؽ5�=�J<�������z�<O-<<����1��<8��=�_���མ��5~����;S���P=}�'=�<<A��m�<�t&�:����Tk<����i= 'Y��3�O��5�=zBֻ~���?��=��#�~P�yɼ<"ƽ�u��� �=|L-��+��g<<(#8<���+�=���z2���ܼtн��ũ��&ڽӇ=�K��������� #d�y>���4=��۽2���f�w�<|*;Ў��J���7"<�D�+=�`������������@�|~?y�9�?��Z�gW$?�h/��ۻ>��N?���>�S?�tO>�P��4:>O��|���v-�]��>��:?�U�R�;?�@-}�>	��g��������>��f?���>k����Z�e�
�✳�8�O��;G��><PԿ�R�> =�8�n.N?c�V��� U-�!���W�ߏ���b =��A?ob��Ä�?K=~[?��e���?����'�o����=�c/?Z{�=$]9��߾?j�K?�i��!,4?�W%?aY̾�����g{�����U׾=<�>N%\>)?�>��?�Nt?_��������='M������|���??����Œ���X|w�f�����3��v`�Jc⿌�J=ELV>p�>�Iƿ��=�׬�`�˿PN����=NkE���s�}$�>@�t�Ї�����A�q�;�_�z>	?�[�@2?!�9r�>޻s�s`ƾǲ����K>O,��>a�`�*Ι����=$	�Xij?`��ݻ�>�!�<�5�?� ���N�Ze�>�FF�"j��jK>"�5?}��?��z>�!?hpx�\��>���k��=l՝������̿��D�ź*>��3?!ޫ�k �/��cQ(?xd>&��&�u�ּ	=�F,���?E�>�(c��=3�g���� ��.���Ѿ��&?/�=xlݾG�C��վg�=piǿ�}2?U���g\�;+"�� J�:�v>Z�>[5?*�����ҿF묾��?�����x�E��>�落}�B��p�=��x?����$N��gr��ɾ>p6�֯��V��>��?�F>�Ux>	��$�k?]C`?ٓ���=L���_?�?�>U����>�=��,I��}�?��?ά�?�ݸ?:�?���n���k��F��?>��"?�Ҿ>޻
?��~d�WS����?8 彑Y0��%?��?�j>?9�@�о��h^V�̋�?�u����a?a��Ǭ�>}(?��G>v�R?<,�x��j�>�/��`?2�p�-��>
n�?G
����X���KW?���y�=($�3��Y�ɼȱ �+z�?�h��W8������Fێ?�������˯��G5[>���Q?�>6��?�P>�n�>Ti��%��>9�n?�����J2�b���Խ�9�=�"��B~ʾT�J�M(������{���������C�?0������hM?��?jc �E�	@)�ҽZg�=�B>G�d?����ţ�?N�w>eP��8�=?Kv�>(Z�=��h���b>����&?�-@>/���ẃ?�OP��1$��x����&��A�>(�?�G��@����?�w��U�4?�)^��g"=Sox����>��п��=�m?��> �?�F��;'r���=!�¿LS?��#�= �����}>�g&��z���׾s;?�Fk;B(��p��y?
I�b7J��+��s�T>��\s?��7�ӧ��� ��MC���w�%1�Q�
��#?��=��J?��^���C?���&���/P<p��� �������𲙽���=��=L��<xz@��Z�RU�<ja=�*<��E�:�=5m��J�=��ܽwu�=Xs�=�%�<��O>�L�=3���T�.�=�M�={����=���cn�<1�ɽȻɼ��k=�|�;l==p�<����¦���#<@�;�m>��>�SJ=�]��z<C{o��Ɯ�ݳ��Pꤽ�̺�d� =�2[<���45�=���;���C��t��<Ïm=����@���@½"Ζ��F"��:˼��(>@ -=�k��I	C�M8���'n��	��_�Խ�޾���"����=�鈽����BPi������O��=qp��M�Ժ�ڏ��1�<i^�d�9������<`=���=+۽��=j����w	�6�!=����z[�V|.�U���9�=޻<6��XH�:j�=b8����>d=��(���$�l<Һ���}=交=<\�=*�L����� \=�%��}J��W��wʼb.�.�5��?Kܹ�W?���K�>62t��K��V��>Ɇ?�b'���>2x�>[,��m�>dNH�����E���Q�#;>ȷA��޿&�վf��<Ѽ������g?�
3>�T8>��I���2�:����`��=h>��:�־���=��&�����T��x఼�+�=U{����?�[��&D��)���پL����Q�>ݝ�ؾ�= �C�%�a=AS?6ӷ��U��: >ٕ,>�$�=h4��|��Mxf=&���˿�����>Fj?Eh}?����L���)x>&9�<.�&��E+>P(?8�<?�ئ>x�5<ʄR?/��?�c���<F>!�?��5U�I���QN"��ۖ?�>�J�<���a��|Q?�c�>sԉ�M~?��A�¾��'Jпl0���\="|��|����?�U��K3>�1��c�&��<��׿���m�֪��Y&�ǥ���#?���0�G���ܽ��:�L���%�?-�r?-��>��᾿��?�V�o$Ƚg��) ?��B�5!>����d婽�}�`�\�sO%�T`[�r�"�;�����>�౾\�?��h?�R;����>>�Z� �Ͽ�xC=��>�#3��Ľ�-�t���FLN�1��>�
=�b��l�����ύ��0����-<	�4o�㙥���𪆽�5��	�ɾ�Ë<ڼ1�Zڐ��c�<Z3�өѽaf>5�9ع3�B
���7���բ�oo��dL�0	�>h�U� z>�G�����탽�wc������ ?x���M�?̰�N����y�ѻ�=���>���Y�>�8� >����I`"�S�?6��K�?%<�=
�켂��>�U,�=:���O�P�о[u����?.�ڿ�۶?���=�d�����j�?<�>�	ſݙ��'(>%�&?������b=�����Oſ���P ]�˳=�NE��!��K.�@	R����2>���ӿ�	���	��գ�Ĵ?R���&�G��賾��ĿB�B���־����<�G�Կ��U���K�ſ��[Q'�\la?�<۽G�Ͽ���<�d��.n/=з��ޯ��H��?��z>�6L�Tс>=�	>#{?V����V�'䅾l�c�'X/�Riۿ'S�i�C=)���*?���R鿊�D�=����e�%�h����>��?��f?��=�en���A���	�Cs�c��>�ff?-�e>�8W?�[��L���k?O7!�i�����L~��_����N���Tf?�V������R?�ÿw�f�Ӄ��@�V?(Ɋ?R�l>�>��*�FsT�q �>�1�����7�>	R>h�>ځ1������>��&%��mB3>z4�=	�=[ň���Ǿ����A3�@L�����q�Ϳ7�1>�ZſL&�>\7U�����u�����.����9�.���>�h�?*�н2�F?�A�=�-s�L�5��:�>W��?��X��bqͿ���?���6�����n��˖=��ξ�x��A�>�.�T�9�</�����>e�>ȴ�=K+B�tUĿ6�y?ˁ��+���@�޽2��(]�>�=R�=*%���<��'�=�	t�8=��Q�*����_����O�� �o�?��?0u���|ҿcbH���?��E����<��p��d뽞9\����>G���'��q�+2&�0}<w���'���I[� L"�K�ֽ�5���%?��7=���=�����Zh�XCl���8=lh?Dn���#�?{\	?��ӽ�A �`�X?�ј=y
�>ۂf>����? �[��ͽ�a�>q�G?�+�=z��=1:�� ;O�z������8�=����ｺ����<�:ؽvJ�>w�h���}��|�����~�?�\�����ç?�k��kK���~ �?�W�>F8�!��`ԍ���?�)�>JɁ��Ƃ���s����`��@F>D~-?��H!��ny ��*��p�[�bf⽀�A=ۦ���?����e��v>�̠�/�1R�>�4��9��>m}�=�I�����9t���T?��?��},�;�d?�>=ş����?E)>�Ӱ���!�=���>��N������?�>aY>��F�^0�>�Ԋ�)KǾ��|��Q�TzI>:�?�5����>Yg���!�H��?�r�?ޓ�~��?t�?�z�Nr�CW�?�t/�l_��2�������M��^=f�����=�Wo<A��
ZW�L�����Gl��!����!��Q?K����>�J徃'&?m>u�Z��`�<1>ڀտ=XF?_d�>m�l�ܾu����=��a?����u? jϾl⋿T����~<�_:�"}��6��\���4�>U��p�>�4�����h��>���m�?
�ýZ%�̟��[��?>l?�+�����ľ�T�����ȕ��WG�8<����J>@M�<1d�="e���=��t�j����Dv�lxr>6-�?x�ž��=q�?�l�4��?�f>a[?i"�?Iݓ���^�L�t��EG=i���q��M�5�E�����J�#V������ܽ�F����+�?8\v��󣽉6><9���)����V?�O��RH2=�� ?Α���=o@�|G׿O!��}0v>Fb�>�|K�Bl?�O�=˄V?�˹��k�>�OZ?�I��ha���@�Vq?��H������ݾ�
���F��;��%��>��-> �J�dvݾpn��x��>@�e=3y/>�Y���n��[��=Rm���t�=C}%�V�����>����k�>0?������OO,�������=���?e����½���Y����9���?�2R?[��>Do�=�j쾲����Ծ���>�d?uf�>���>r�>��ӿK��=NG>�?R־M�}��f�=�Z">$F�>Uz�>,_�=�M�>F�G?x������jy?+�w?^1?,rѾ�*�>���<dr!��/�>Y����Q��9��qE�����'��\�����|�<y��H��~$}������?lM��Ӭݾ���?�[v?���=��ƿ^��sᔿ�a>�3��X��g�������<p�w=��=P�3�E�<�=���'�9�����M(��N�����:�������<�fؽnf�<�7�� �D��< ّ<+>Y�d�$����������':���<�z�\��=w��=����=O�Ѽ�ߋ�L����J�[����5�������"޼`_�;���7զ����=`<��Q=��u*��[��,5=��&�^��<PkL���<��g�*,�=��^=�|Ͻ�q��7�\��ZR���2��6�=��f���*?\:�u��=�����W�>�5��l��D�>}��>8E+���>�F(>�v��Zf_>�H���wK���پ9�(�L�>*�x���?>��5�\��v�7>t�=���O�ƿ�>-���O?���)�>7��<Q�=�>޿�ы�
�~=�1j��g.�S|N>r���3�M
���ļ? ���h���0���ξ�����P?�h]���m\I?�d&>�h��?l{	�Ns�7���,�ĩ����?�=����=/�L=���=GH@=�m�<�Oݽ�5ƽ�}=,H+�� ��p��xʽ`Oӽ���=[���g��w��P �� d�c�P;�c���˱=�y�N</��h�|�ʽ_Խ�(�=x>o=���*ӽ��<�D:a�q=|�S=Q�i��Nb=��|=H��Hb����=x Ӽ���<��d=�"�ː<7W�;�A"���z�� "I=�~=�@ڽ�-�������Ė��[=H(���:��D��6V=����V�p=֎�K��=�����+���龏��=;�����ž��?M�����������2 �_��>í:�$V�>J�A�p01�fI)=!�˿��U�;�.?��`dM=i۾Q2����>r�>�`�P��)F�!�ο������D�dv��v�P�x����W��̅��~}�o�=T���ۦ�x�>�T&�x4=;����)Ӿl�>�:�� [�P�c��z9��$>?�>��.7g����?�6��nQ�y�M�5	��o>�����\�=��!=��7?Ŝ=�*��I+F>��-@zU�6�j����b�꿙�r��Օ>�ɴ��̀���?�؈=�A�,ݳ<�!��C�����H?!�8?� x��#?PMG��R���j�#��?�E�>t��MU?{yʽ��<������M?�{v�8�0�)�>G!,���I=�@�|h>;1⾜�E���龼�D��9R?�y��q�W�?8�?v��ظ�?�d�p�<� �lz?v[%�T�
>ɬ���j>�45��ln?ǇI=�m�>O�@h5�?8�>F�žPē��C����쿡��>��ơ|�夎> ��>�x?!z�=׆����?�x%��7ӽ�(�=�H,?T�B�[�����\?�-@�v���=a2��9�:?�����>	
�����>�v@�NǗ���������L��ws>N��=V���]�y�7^@T��=�����b��Ö>���)K�?��V?�Ա>���y��?���^AW@P�>�?���>U�
�e��?�aM�<�?0�=�B�;@k�`�+=h����V�3���c��
�="]�:��M������罶����Qh��勽씶� M:�K���ս�XQ=ե��Q�y�༽"���������E7=M\�<�C����=oG��~����2��4�m�(н�ؽdqX=cn��m�u�=�λ<��,<RϽ0주�'=1�q=s��<t�f=���=����9��=���X��=EQ=pk�<�_���$�<��<���=����8=R���������E��(��=���������>����(>\ы>ɾX�����<�k��k+�����<�j����P�VN����=��X��CY�=0�����<�O�����>�?(?*��#��q|m�Go⽄���D ����>s�x��I�T1p�q`ýcR�`Ԁ�6b�������>��
<�����i	*��>� >tZN>嬸�> #�d+	�(�ܽdR2?��w��ӿ�\����.<v�;�%)۾\=8�O=:Lf?/�%?}P�>�<� 6=�U]?� C�c��Ẹ�߾�c���վ�������>"8�1��?�'?�ś>��;?�I�=�d�>�t��)ۿ�?�9���v?�T�?j�?	=�����E������N�)\�?����V�?���=V��?馾�L�������?��Z>a�?'����>�¿=�-?
ۗ��W>W��P���/�?���?tQ=���>�l���my?�\?&���l:�/��?j!)�:��<��������ԫ=P��<����@�ѻ�U�<�@��@Q�;fJ�����=����H��NF,��뺼 ��
f��W~��`�=�c���>�=�Lн����<�s	���=`:� h�;(�A�06-��:���o��z,�=.7�{�� j.����Ro{=����d齀�#��Uk:�Vg��ʧ���[�Zp7����=�T� ?ۺ#��eW�Еѽ7���
�=2-���
�;S
�:�@��㽆U-�n�y=ܘ�龼@�+>������=	��>̾蓃�#1��˿�w�>�;��)&��h�>�)?(cR���><�(���2E�=;��1�=��s>;���O���R>�Ҷ?�=���Me��?�a>MT)?�Z����0?��1?/��4�#�"��>p8�g�`�Z��<1S=��=�K���9���?���&��&�>}��*�)�蘨���B��n7?C��>W@���=p��?������ ��<ej��m���,?)$}���ͼ:{5�U�<�`M=g���ǽ��<��������Zu��8�=�xZ=c�sc)>���!���!~ڽ��=��7�F�Z=�U��(ｴ��#]����"�ݹ�j�<-.2��x��9>�ɖ�k�?���/�p%���@�=v$�|:Ƚ`�_�P�轌�=h��<<�r��6<�O����=�O�J�r�S�:=$� ��%��g���<��u�&�	� %i=������<����[T�j���U�^��=z2$�kJ�=`
�5�g?$/>�>���4,�>��/�;�E����>�zž�庾���>p1�=�9Ǿ��Y>JR��(]�׾��Vʊ>��?>�F¿^�>�O�>?�L>)[�>�gǿ�[��i?��o?�F?��s����>4����<��}νV�'��ṿl5����<dԽ=��ҿ��¿.{M>�-P=��!�+�Ps�У�-�2>8�>����l��>d!��sK=B�3=��k�o��4�þ)~�<�%���Q���/� (<�v����;��˄(=��`�Ajy<�N��-�伎_r=h��B0=iW>^�"��Ǔ�{�2=��9�]���=���=�:��s��kZ�g_�=7D���̼���=�36="wŽ����˽�7��è���N��:��P���3f=���g�����=�aa="l��!� 9���΢=O�1��MR��Cf�[d	=ol��@^=��=�FؼN�>��Ž��-=���;��?=�坽�����;�]�<n�-���?���=�?�N>�oξ�==J����>#�`�������>ѭ?=����>�q࿝�3?y�i� p�_=t1���IG�?C�|3U=�W˾�?�7�K�>�pV?*B??������� ,�n@s>��;��tI������0-�"�ʿ�.��ȷ�<{�߽(k�=R�?�5�=1S���ksC�,�"�ō��ؿ������]�l,�=��k=�ǿhۿ��X��4����?6�?n�'�m<>7*==���>��>пڿ��s?���d�>���P�>0��<�Sսz^M>,SB��޾|+�Mg?�>P0�>�Ż�i���La:�?M៿�׬�I�`M�;�g&�.��=�Ѿ�y�>��l?ц>&o���Ɍ�g=ɜ�� ����=�; �T�����"�=�Jn��?=a��=�0�=}a�����@�>Y��������=->��)�����]�=%�?˦`�����4}�������>�1�����)����<2�m�Ko=B&
�`I<�)�^xC���ɽ@(���%���I�={��3�½�>�<{10;�Y=թ��W�|{���->��=�}�4�����׏ܽ�Q�� �y�5������H������u�����靽�\=i=�����=[�����;�=ʈȽ�W��Z��E<����=}^=���K^�eAP�	ǘ��;+A$���º�8I��=?��<<�_�<\_�� �����=
��<؊�t����Ȧ��($?������ ?r*��s�$ʿ�^�[+ ?�M
�Z!�y`C>�t;?�蝾���>���5eK�p�����T����=��4��{���Θ�����A��YB�Y�!>y�(�ʳ?�'A>~X0?ub�V~?�!&�������<����I}��P�R稽��D�7�N:@5Ͻ�T��0��D�1>|��,�t���X�L8��IU�>,��=׷�>��_��=�?�I+>y���<�4$}=����c���Y??�KT?��1>g�I��&>�����=���>�?��s�wL�>
C�>
]���];>�x]�\AN?����y�E����=�����??�ὦ��=6�[?z
������j ��c�?u'~?HG���8��<>x��s7οk���m�j����ް��c?:��=%�F�����sT�N��=Ӯ#�+l��p:? �f�i?6���d�=U(ʿ�I�F�=�W��M�?����ae?�=?ℿ�8����Ѿ�j�Ph�>F�����e��>���vo-�4?�~��XI�=QI���=��!*=/���l�ۿ���=V�?<�ƽD�f�Qy:�1�=Rar��{��c������i�$��y���T?��>���>{��=4�e���=���X���	����?�"�=�}��`
���->����G��'x,�8O>���=p��=5���n?�,?�i�?��տ�s?�5���?�=X�� �y��x3�t���8��� ����?��K>2����6���"�"���<G��z�J���4)��oP=�~����M>b�%>뾰���X=��<�=�=8�W�>�W��о1>�>Rҽ��<�;�	�x���L=��=����e��̀�p�x>pI����<'E�v1�=�9;�鎽�^?<	醽���)���=��{=p<W�/���<=��r=������9�ڽ˓�V��dN�<�,�ɌM=�I�=�wg=�P�����=tü	��=�l$�򨜽A�쁂=5�5�=��>JҠ?E)�>-��X�L?&x�t+�����|�>"�
@l5>�� ��b����>��>ʴȿ�I����?�� ������>����䐿����t�>�u�mu�>�E�>�[9��6��*=��s��a�Q�$�^�??���ن_�K��ac?�5�=�:!��8?�;�W?~@��n#>k��>��V��u>d|�����c_�i�>��r��8����1?��W��wT->�����?���4��{��aؽ�=a���9���^7ǽU��Ba�;9����.��n�={�Խ������]��H��v����
=������<8�E=�����q=ɸg�=^��O�9����T=I:��5G=�3��D��[�� �s:u�+��<�D&=�G]�1�ϼ`:\�0�*��ۥ=��H�j�=��=�=I_=��
���s��G�nRs�5�νm=���b]�=_3�����v;�������"�6������`;Rb���e>���<�4�;�c7��ܯ�����7�����=��=�w�==Q�J�~�`�����=�u����=�`@��J�N[=v�=��
���4�)�k��Nc����6=��ѾP��<�ڎ�V�A�%�=͗�������Y��&*��dX���'�����Q����/W=����"�(�_e#��ڽ������J�8�$��w/�cz�= ��?6Ƽ��#���[=Z�����>^�-�^Û�,~�;h�<F��=cb�;2%�����?8�?�5���C�wJ�EA����6<���ʋ0�O'<"Yм{A2=�=�=(�b���.�2��=�Af��4�=�_�<��#�G78��1��`Q��}K�n?^��=|=����ջ�r� ����)�kʼ���=�$=N�j��ܞ�Y�P<`�N�2��W���>����=ɟB��O=u �=s����Vn=YWz��r1��;t>�����������d��=�O�='�A��6]��c*=M�ټoh=P�弄T�c�+�`�P�=&S�=P��=�)�5����~�<A��<�<=��#����Q6]�q4�rр���������ļ����n��}������>l�=�A��Y1���<��⽰�μp �=�S�=ġ`=��;�5��0(��[��g��&��=Vk>�BP"��	�8�D�L��e�^�M=��̂��=?Rw����Y���d��������w���0��,���آ=���=Y�5<�_��!�"��
:���=,��=�+q��$���=��p�<D9=d:<�4�c�w�������!�}=�x�=ˌ�m�<���<D}�W�.=8�m;S��;-�<��=3�<�IUW<�! �f��=�&#<�����< k�=���<�ܽ��q�(\=?���
��o�M��P�X=����\5���<p���ݣ����<�<�=�"�=۪�5ӽx�B��'*�U�=I��=%�!�bᵽYN����;# �=�T�<�g�=��E��<H�J=:z�i�;
��%�@;�*?cd?p��<.^o�tvW�Lee���Ͼ17���c�>8z�>�kU�-'�=�D�=�a�=�9>)�2?���.�?����~���KZ�v$
����>�i_��w�>��~?/���
n�E��z�?,��[l_��n.�&ʉ�*X�?�v��U���t>jL�h����{,�(��' �?����n����+?{�'���a��ԛ�Z�@��h>�fǿr�?~��=$��z�>�M��t��Y�~�="�P�0�
>0�<GP~=24�"�%�2D�=��%�Ұ����"��a6��7�=�=�g����)��Pɻ,�������?ѷ�v��[�9�T�������Q�ڽ����~�9g�=y���V�<dre=K�C<z��< �潾�(��� �<�o�/���C�=9ԡ�Qt콍d�С����4<
Uн=���ڂ�y�=�3���Y�����S�=x���;�;h~Ӽ�_!��{$=CuཬQw��BR���4�g���+M=ڽ<��|�X�C=������F�=_��= ��!��=�b��E��۽��G�=V(y�}�=|���Oν�E�=A�Z=�"����/����=׼�?��5�=�e�<�z�<F�`=�]�1��\�8�g��(/x��'-=�_����ZA��e�<{��<D�׽X���O�^�W��m���R�+｡�	=��=p�=N�<5���@z�I���Ì��A�"�Ma��p����=h;�=��g<ۦ���Ƚ�^��+S�ᤞ����=@~=�T�=gZW=Љ����޾��>�����s龰0�� !?�ؑ�E�<�r4>���> Ih��	>��y��R8?�Ȣ�� �I_>t�s��P?}�¾��<>�A��p��l@'>C�;����>fݽ?{Ұ�����M��?��oKz��s?���W,<�xW�2O�<�ۦ�� $=Ԕ��N\f�dt�=����&�����J��pZ�><�L>�_h�˫�����=OM>y#H?�J�%/.><�W���>��4�� ��Hc`� ���.�@�N� ?_䳾���>3����e>�)��K��nC��}2�?�1�о{ߤ>�ǻ���>���=6�Q�ғ�Y�4�N�1<%4��f־�����$�� Z=��>�z�>�*����ſ���!=�>�ǿ-�6�`㞼K <_�����W�Y���R������ ;�Z, �����*R?~n��&b� B�<���W�$��>�?�ϱ�՟��Nؿ�)�����>4ċ��!�=�c�>�m��*=?�����n���M�����=X‽�'�=��ٽ�9�m
�T=$���0���X(=����@�<�I����=J�E�'��_O<_�����_���︽_=��'
"<����OX��䲽�g�=@
�=x�=�NA����W�8�=v��~�����۽װ���Y�n���4��=�r\���ĺ ��9�̛;��Ͻ{���1<�7	=$��<�W�gҼ��9}�^)�=�7��	P�=�{�Ja=~ZS��!�ȸ=n`�������>i��7��>JkD�o�?HF�妌�32>2��>��'�^��>��n>-�����>>G��sW�m"�=����6�=��)�)Ae��)�>�N��8��
1��ؿ�r ��%>E�?LQ�����>���Z�AJ�:_)��〼���v�>B_�>`j��\S?\����N>�'�=��翺� ���/����fO����g�Ƹ��"+���X@�؝�����$>��,>I}�zO@>|��>�V'����>�t[��
F��?�0��=�@�=����f=S��	�i��v�u=��m=V��[o���;�+��=bh��ӓ�a'��V;�b�h4����
�$���+���x_=* ռ���=}d�$:�����y+���
��g�=T1ս�'=N�����@�иr=
��KoZ�D��#�!��sD=D#,��	��� =`�=$�<��<γ#�|b.=;�;=�A ;�끽B���=��?���ѽ�ԛ��ʼ��;+<��J��4�����>�ʆ?40��J�T���V?�#�=�@=o��>kL?'�`���i>��>��S=�Q�>�0v��zE�����>�����@>�Y��f-���%1n�j���'��>��}9��tM?آ�=?�O ��ꤿ���=����W?:�~���	��W�:���2��=��!?�]��?E�=�G������7��X��c>1�����̾2zA�d�ҾT�;m��>Q�翚uV>;i�>�@־�$[=^V0����� ����H��R���������H�<��
���s �=\;�=TY�Ij�= �8��콀�n;���<��Mȝ=����?�=�U���]=ݯ?��J����� �2�0��Y��~`���ِ=�����׽�6I��r�= Ь�'{ӽL�=�<&;,��;�ϼ���=6�%�4�������"������`�i=;�=�ƽ��v��n�F�4�L�#�����ڽ�2<P�-<���=�x9=��=H>	�:�Ƚ���IL�<�zj>e�Z?�]/?	�>��U���4�p0>�OA����?	��>�y��R�>]=�>ۈ��WՆ>��&?��?����o9�z�>֌���ڿ���r�R�]�?i[�=��¿
�>��>�#�?��?Ҕ�?;@�1r=�o޿�>��.=I�5�zL�`)Q=D�?�/>��=`�<V�G�U��=-ɕ�g����ÿBm�?�n��I.޾��@-�>a��?�G?+:?���?aC)?E�O0i>�-a�oT��a��ӎ@�*{?)�?
Vo�L���?��H��>�F�?0L���َ>�<?(?$���@>��/8���=l��>ӕ��֜;>��19���k@�+l?"�^?|�׿Nu�>l���@{�?�6?�m@WW6?<n������2<5���=r]��}Ҍ���@���B����� KĿ���_*��dM�������e��eg�?�k��x-?i9?�k��|�۾]?�T��4�i��>�S��i�>s[A?�ӭ����<@���S�>�>����$5�3�>��e�P=�=>�`;xac����>Ņr>L_/?�5?P�"?�Ov��^�>��<n{?쮔�]�W��B>����Z��j��0s���Q��?3\��¿�	'�*���WB��E�ʾ��=l�s��Z��G:� ��<})����a�T��>D@�Yk�������=�۠����/���^=@�<>�L���<A+�?� b�&ۀ��7��"��/~>]Pľ�F��E��������?� ظ?6ɩ����?П��D�=>ɘ?R��>��)��s�>��x�D�>��?��@Qq?M�l��=�r�}�?�5�?;�>��k�?�"�e�ʿ�� � q�?�ظ?�Y@YH�>Z�?��̿��=�ؙ�̦=�
u?�ٌ��E@`ཪ珿d�c�X��>�����3K���.?�f��!f��O�%@��@&3y?�$�?;i�?p,G�A��P�,?+�̾�@�YO?���R͠?C��)�}��ۿ@�#���A�D�??��ž� �2�a�ȷ���.>B?�>��#���j=��;?��x�e?M@��_�d��������_�<5O� {s�/e��_V�B�����C�]h����?^��>Ͽ�Z�>񵛿Ӕ��bU?���J=��J��6�?7r�Q���PU����?ݒ��(��R��=X噿�d�.J=�� �P
W?G	�?'��<��{?|��>@�l=�Ͽs��b�<��@�����>Æ?ٍ?d˽��6�l{�>;���ى�>��p>������.>�$��e���]�"P�>"
r>.�<>�6���������Pd?z��<��'>��W>�х�a#��E��'ޱ>�*�7j�>��	��୿ �>p=%�ڽ��.��M���R����=�a��<�n��Մ>!�2�>Ǳ=��>�>Q�M
V��O�<�\���>���>^����>��<?ȿ�?�?=���$3U=�3?��l�1���?\����+�<����!��m�=f+�����=�~�<k�n�0��*o�7�����?�zZM����;������<+J���-�J�/�)=����#˽�8j=u���h�=\�<�=���(�%��lm= 9P:�c콄�=�0�=t���L=��=��������@��b��V��#��\4�=_S�=\���O��p��=�q$�=c������mﻑ�����������k��w��������i��	��+��2���_���؝�=���Q"<|⑽����?9<͹�$����侎����,��R5c=߬�=+�>Oׯ�Fݓ��4,�5�A�h�㽊.�M\9�**"�²L���㽶81>��SI�ݯ������'�$������<E�=�	��Jr6��h��������ڽ�*&�s�̿ �:؇";�5�>)�� Ȑ�[^w>�g;��WмZ*�r���c���EK���'꥾�B����=�T��L:�༥�od?��z���m=Ʉ�>�vս$�?=@Hо��Ҽ3��|��A�?�Q�����>�o/>A3=w
>��q�:��> JU?���>A��="�0?#��9��>;�[>����(Ų=�v@��~=�aɾ���n��!Ӿ�e����=��-��w|��%�;O�?������� l�4���Hy��A#?CM�����=���>�����B���ÿ;����w<�Ig�wf;���!����{�h�bR]���Q�eѾww�<��lfk?.�������� ?7�S���>�+?�(^���<@x4�f�:�ƌ!>���?�O�ZK.��Ͼ+�`���@��䝿���t�=l� ���ѽ�-��D���e�8>_��<?��<R��h_��E�8�
��a��_�����վ.���Ą>*j�>0�T���ɾlٕ=��>��=�k�����ѽ$?�H ?��ֻ�C?�x���?@�9;ے=�u���.�h>�, >�#�[���ul�:<�ʎ�=@��=<���x�L��=N����ƞ�h�����=�落4�*�bz3�r<�=`M����<X�<�u�MŽ�v=-D�o��2��.<��=�I
���z=�%=99D<��x�1�thy���=|�x�l�콱`8�[׽4�ܼip=����b��`��;?m�;]�=��u��TɽU<�����$�<�W��8G׼d�2=�0�r���~="4���Ъ��~*���(��4�b��^�9�Q�\=�j�����B��47�k��<����D=?�!�A�����6L@���<��>�ј�?9?���>Y��?���d�,�[�S�}1�>~��?l ��<�>��?0�j?�w=փ)>A�>�м���K�>�����-=���?#I��?(_�0-?��+?nʹ?�%�?/�B?�,�>��©��`ʾ�Ͽ�X�T�>gQ�=�+@��=�J�?O�i�E�>�#=�C����>����?4�[?Nk�> ?96��7�?�f�<�!n����vl�\��>r��?<SV�;S?�]��-ҽ
>�>�@�8�?[��eI?�)>y�\�K����k�}H/��t�>��?ʘ¾��!?�򿔲?F[5��W�`Q�=����^6�����>��R�=3��F�BkY���쿯���*�8�辌���ڽ7}�� {�=����	�o� �=Z"P�M����p��hvp�"Wb���.?��>�E=��m�T?��;��v�m�`�/>�q���,������.޽'��=)ܜ����;�� �=AM�?�ӈ��ʮ?)�=T{'����<P5D=ђ�=��M�J���Т*� � �e�ὒ��Y/�<aD<���<��ڼ��=�������<�d���r�<*'�=e
%��$(��=&(�4�Z�s��ǽ����曻�7[	>�,=���\��X`�=��˽Aؽ��2�V�7`~��y�؍	�nl<��j��GB���M�=S��2!Ͻÿ�;O�=ֱ��I2=�4������w>U=���I� ���n=���B&F����Ւ��	|���=�8�=!%�����5H��ȽB<}��N�>�M��J��CD?�k����[?O�ݼ$�=��?�u�=|��<�j�Ľi��������~~ž�"��}��\|���$?�8*�p𑾛n���L)�K	���i����>7ZϿ�P1=�7q�w��>��(<�N���ҩ��m�hAν���>8Eſ��A=��=Ϸ�����	u��� ��f�q-�?��O��۾��>��(�����$A��%(b�?(F��N���s�?����P���=�н`v���]�<�{M=��<M��<�)�!}�=Y|��E=���ၗ�.�	�E4=<|�=�=�����<���ֆ����n������E3�!�Ͻ7i��;�Ľ����T�<��[=!�޼�y%�j� �@?��n�( �=.�0�@��|a<d�a�W=�=�==yٗ�Qw�=I��\�<C&�<���}nԽ�1��m��$�ԣ5��4ռl�ؽ�@�=���g��_J���ӽ
R�<�ٽ�8��"�'���[��>����*C��-�>�>�U�<m�2�<�ܽn�=����1��#Ŀ��
��a�>�ѿ�	 ?p)���Hu�u�[>�)��i�ֿ?�*���J>����~�4=:�>@����>#�G?v+��+�)>���.z�=�tP���u��I�=(ќ���������c�=�Y�j�� �ڿ8V&=�ގ�̼w=p=׼��'�t�ӽk�V��!��
�ֵ>m|9�RԽ�ȫ�ٵ*�Ƨ�h��=�j��+��<W����͕=��w=[Ή<�6���s�Z��=�Xн��F��;a���!�;���(�P;kl��<;�O����l�=*�V=W@t�F�=�ǭ:�����������ý>)4<*P���͖d<c���ĤW��Oνn��=�m�=`g=��ޅ�<����J�� -���;�8�����j��=�*=����B��������B��<Fk=N0��oz=��h=��#=�:��N�Q��(�q�W��=	_L��C����=;�?��?}i���ď>`� �Od�>m�ξ�j�o��>;���1�`�>P��>�#� ?�>���Xk�>�`�>`!ܿߏ�>}�)?�L�c6�>�H>�+��?��;?m�ܽ??6��Q �>���>D�����U?��==.7����>�>5Z��t�^�۾���=<|?A4*�t��=Y�+�j12�D�D�i霿���?�~���?Z�?u��?!�>�����5��U�,�Cx�>Ȝ��5�>��\�"�����QZ���>�=�0�Ή���ma=�|�I�C�;ݡ�p �T�q�2��>g�?�B1����D���Da�fƩ�uL�ng�?E���y��k'��ϩ���=H���PcϾ/����ݽG�>����7�x�9�ID|���ξ@v�;�����>8�ӾD`.=�
��� =�M#�<����13��%���!�� ¾�w�D�D�֫��!���FI>	A=�c��b�$�9a�=�Ҿ1�6t�>������^p=�����?$
D>�J?��=���+jH�b;7>��?��z��IQ>ܞ�>�I�>FZ�y�>)mT���_?���>0&���k>�ܚ��hp���>�d��Y��6��L�g-�����ύ>���<k��$Uk=�4ҽ(���o0��k>�KY�T�����@���O��>��y�F�> �ֻ�!���Ͼ�p�>����Ñl��a���徯%`�&��q<©�?��ʾ%���t>���>%����҆���!�=I �Վs>Z�?j�=h۔��^���?i�?qɧ>�kp�2ǿ>�Kq�:��>?�=�c�?�z������l?�Y�=~�k�Е����<��пl>o\��f� *���}{�u*,>`�?�"�z?����g>� ����G�>>`����E?~���d쾍�x��0��)r��+�>���j�>�I����>�ݿY?"?st��G�����~�?|�m�ϴ�?Ò�>|��>PR>B�?�A?W���(���ԫ�>���q0?f�eV$���S�8�>ϱd>�'�?���Y=�/l?
v�>Φ�>��+���>}þ�@H��� >��ϿQ$���7���7F���r��j�U>7�!>Rֿ� �>{�>�h_�vl,��f-���5��������V�?>���>SkԿxw�<�_����1��c�?�L�<�����s�=T_�i/� HȾ�V�y����h��M��t�:��R���������=-7���8?2r>��Z��<��>= �� ��< kf<�l�D;�1�5ỽ��u=�x��������<��.;��潴y7=��O<�U �`?t��F�����=`��=ғ�=�}��$�=���S����*�=ؒ=�z8=�x��7�N=�|�y��:�,��{;�2����s�o�h�=�ތ
���=O��<�ཀl����=Pb�<���^/��l�a����@���H=�⿽Q�M=���D���C�Wջ��g�ߩ�4��=��<���; �u���ɽJ���_n�=,�L�/=�x4��[Ƚ\H�H���нL�l<X�ܽ�ZϽ�r���㗼-��=��=�W���U;�!=f��b2l�G��>�e=�a�=�2��HU�����l<PD�=d�=�jҽ�������=x�˽�������}�A=�N�o T�2ؚ=Eu;����ar�8��=��E;v����ƽ�%>�fZ����.�;��&:�#���=A����m��ap4�2��t���Z =�h'�o�\��=j���(��\+`�y�.�%c-�7f�	o?��?bV��G��1�ѿؕ�<�}=U��>y�=�;�nP�=�w��&���R騽@.���ڃ�ɐ��"?_�Ҿܤп4�F>�;��^��$}��y�?�����9?�A����?��+������R2��	�>�!X���=뭱�R<��w-� �9;�f�_�#�C(�p2þH)">	=���
ھ��O>�� @1�N~�ܓ�����?n��̾��>@XT��M�>D�J=*����=�"�=��ҽ͝3�h���^>�ԣ���[�=��<g�ٽ�<�=ނ<Gj+�0<;2U���ѽ�g
���-<��<�����=���P��/���w���`��'�{�˽���=j�.=�����(���=��!=�+<�;�=4js��><�cB<<���=�A=�Lo=(y�('�<����,=�=���:�p0=\ǻL{D�a�	������Ľ����V+��+>�P�<�d��s� ֯�Dv��N����>=���=|�;o��>3�Ҿ�� =��?Jcy�}^��T�5?s���V��!>�����
?;9���!?a���gr^�@��=�ai�H�ɿ,у=)1}>�G_��<�ձ/��\{�? P��⾕��/E>�Ҁ�������5��=BBT������>�T⽁Ȏ����Sա�D���ǅ����/=�ZE� ��>'��>E�&��������� M�=�v]?H��P� ��:��ٌ��G��>����T�qS<4Ё�=�>����k���=��������������>(�P?G�c��A��	�>A+࿗ /��4I��d�>����q����hf>���>���>X;:�������L?�P�?�����P�ܡ=%V|?7�z���;?$�?s�?Ty���1~��D�=Kg�<�O1����=�o�q-P���a��0���3=��a�VQ)�s��>@����"���y=@�#���>���YM�=dv��� ?�M=�N^={�;#!ھ52&���^�PKs��� �   �  PK                      archive/data/3FB  �=�>|=�51���?�7P�<���>�T�=���>:~��}��?�r?v��P�>�罛��>v�����4掽��4�;wY=mӽɮ>G��&��/���u���z�>��g?B�r�qe&�ת�fݽ_�
<�d���������v�>�1׽�+�>����&ս�I?��>ώP�+̻?�����6���H��;51?��<��|DZ>�Q���j�QR��[U>����y��W?a�%A�nc��m�>��Ў� o���<���ɾ$�����:�,t�>�O���y�;���{?���=Szƽ�n>t��?p��&]$��Z,���n���5�WA+�,����C��)����z�5,S���l�?���aC<�aH�2lҽ7�Ƚ��?ƐH?�>}�T�@��?Ñ���#��Bg��c{����H����?AO���l �O����f�;b����%�k����[�=vE���p��Z2#����P'�F;8����Q��>PK��Q�      PK                      archive/data/4FB  k|�=�����Վ=Î�?����n~�`�?h���"�?���%7Z?d�&@Qω������:jο�C�?��<�f�?�2?si!@f�ȼh�ʿ Z��r!;��Ѽ�>����?�`���8N%�X�=W�Ŀ���<0-�;Qռ͈���д?-��?t&@���;�;��̜*?l�"@�@��>����&��=��μ�H?w��?F�[? ���@67��5�)��Ԑ�/��>2�F?�G���<k@\����?�ɿ�C�����j�;���p����0@a�)���O?�8I�),$@�~�?�);=Zn��>�<?�t�=�@@=*;z�m��V�*5���堽���命\��<;E�?�)��8"=O����߼���P>u�<Uߞ�?*�?���?��~?\@���*�S=2�h�2���P?x"�<��U?��L�ą�:���<�����C~�G��3)?g�&�k���͙��:�<:9�ERּ#˾?��ῧ�v��"[ռm��;����<<d]=䅘�m�ʿ������8?�b���_��p��ݸ<7�b<p����={Ͻ��?Z�u?�[O�!@o��<F3,=��K��e����>�:�>���ȯ;OoG��ؿ���<xH�?�1z��j?��@?VѰ?A�O>4U<�]����>��;�6�п��>��翉�@Ա'���H��mM?�A�?��?O�h<[KP?�*ſ_?ҿ��?�m?Cd����R�1���w���b�B;���?f�g!ÿe���;��?��?�;�c��>י��
���� Y="CB�Q���ʵ����?�p?�'8?�U�=��Y���Y�>*�=]�m� b<?]��� ��D�z1=�������?��Q=�|��﮼�i�m��=������<,?�Q?z��?孆>�X^:�?6ێ>��?�V=�C?��J���,��1�=[z��>�z�;R�e?1{1?b��?b��?\?ia���EA�q%���I�>L?�ſ�G�X�]<�}�<h`�?&i�?�&�����B��?��v?���?���>����
?�>�:?�����?�����d<A�@��?*������:��@�׆<@��Q`=��D?�jQ��j��Ps�����=t,a�J�����=�K�$ �7Ԃ��G����ؿ�G�?o(��h!=K�*?kl����R^r?���~��
䳹��Ϻ�N(?�ɪ?�ӱ:@L��?؞`@�&ݿ+1?��d��-�?�����)���)=���?>n=��^?���ֿ8����5�`1ſ��]������O982>��!��\�>k�H����=��ݾ�Z?K�?�;}k���y�;�<'g�<���'k��A��t_�����;�Q?��+?�-=���?r�4<B���,K�b�׽n��>ƴ��si?��&@��@q����?�B�??D��[�<렀?��5�ɻ7�@]�ʰ�?�_���=��?}���߿o+��s=Y/���p���3�R7����<!�?���M<�>�<荿b�?��=Q�1���@W @Fa%�ZA�=�74�g��?��?�Iq����?'�%���<;1@�W���H�?��;}��?��<�l<��kA����>�@ Ռ>����(�<�@<ә'@��D<Fﾢ@�o�@��*?a?`�ث%��A�<4י:0�?�@*慿���=�><��D@�A�^v%<�>�C�?��¾5�R@���?W$@��>��ѿ�(@��;�e^����>�=�ߤ�h����1�?�T�����3=~�l=��п��m���{�	1�?��<Mk@���>�w�����?����n��=�=���=�}�=�'���!+����z�ٿ������U�T!?���L���v��?����?���=����?ň���? ��?�,@�i�<��� ��?�}��q$<��?��@�i�<�ĿI�#��Q�?7�ڻ�H��S�?��;��a��?̮����<���?n��=� ��Y�?PKNh2�      PK                      archive/data/5FB  a��?��?e��?!�?PK��      PK                     3 archive/versionFB/ ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ3
PKўgU      PK          �od�p  p                   archive/data.pklPK          7�C�                   �  archive/data/0PK          p��b                     archive/data/1PK          s��� �   �               P  archive/data/2PK          ��Q�                   ��  archive/data/3PK          Nh2�                   Ж  archive/data/4PK          ��                   �  archive/data/5PK          ўgU                   `�  archive/versionPK,       -                       �      ҟ      PK    ��         PK      �  ҟ    