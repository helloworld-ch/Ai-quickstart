PK                      archive/data.pklFB ZZZZZZZZZZZZZZ�ccollections
OrderedDict
q )Rq(X   conv1.weightqctorch._utils
_rebuild_tensor_v2
q((X   storageqctorch
FloatStorage
qX   0qX   cpuqM $tqQK (K@KKKtq	(K�K	KKtq
�h )RqtqRqX
   conv1.biasqh((hhX   1qhK@tqQK K@�qK�q�h )RqtqRqX
   bn1.weightqh((hhX   2qhK@tqQK K@�qK�q�h )RqtqRqX   bn1.biasqh((hhX   3qhK@tq QK K@�q!K�q"�h )Rq#tq$Rq%X   bn1.running_meanq&h((hhX   4q'hK@tq(QK K@�q)K�q*�h )Rq+tq,Rq-X   bn1.running_varq.h((hhX   5q/hK@tq0QK K@�q1K�q2�h )Rq3tq4Rq5X   bn1.num_batches_trackedq6h((hctorch
LongStorage
q7X   6q8hKtq9QK ))�h )Rq:tq;Rq<X
   fc1.weightq=h((hhX   7q>hJ   tq?QK K�M �q@M K�qA�h )RqBtqCRqDX   fc1.biasqEh((hhX   8qFhK�tqGQK K��qHK�qI�h )RqJtqKRqLX
   out.weightqMh((hhX   9qNhM tqOQK KK��qPK�K�qQ�h )RqRtqSRqTX   out.biasqUh((hhX   10qVhKtqWQK K�qXK�qY�h )RqZtq[Rq\u}q]X	   _metadataq^h )Rq_(X    q`}qaX   versionqbKsX   conv1qc}qdhbKsX   bn1qe}qfhbKsX   fc1qg}qhhbKsX   outqi}qjhbKsusb.PK����    PK                     B archive/data/0FB> ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZYw�$[?q]p�zN"���E@��Ͼ�	�=*��G ¾=0뾜� ?S�����/� rE@ɧ����=�z�b�������>{g��B���+E@���KG>$�)�c�������>!�'�@n�z�B@3�ۗ >�n$�j���}>ھ�%�>��d�gP�l?@�ȾR��=�����㾍}پ��?�(��#�j�A@��ɾ3�7>6���]��N۾��>'f�BJ��A@Ld���Q>^���޾}������>�bP���+�F�>@ty��],>��wN�����M��>�3����wC@�s��i�=�&�K���x���>w�|�կ�&�F@�ƾ��<>TS!�}�����q��>Wܣ��>"�*�C@,�ھ�&>>/���Q����>&�$�1�Z�C@"=���ˤ=�����-�ݾW��>X���@� �E@�j���M|=F��)ӱ�Iy޾]`�>�c��b�)��@@�d���_I>�/�]-Ǿ��۾�A�>2i��0��>@uJ�!��=�u��׾-?	����>��T�?���F@o��^�=0'��P��.�3?Rҽ��]>릣>���o�>��?�񣿎����?��#X>3��>���y�	>��?^ ���i��&�'?�J	��̠>K9�>���;�">��?X��� =��H�?ʄ�Ha6>���>���ctL=w��?����.�迲�4?�b%��
>>k$�>n��em=Qb�?�L��*�?f�V}�>��>��#�=���?J���8
�x�(?&�#�4�>oq�>0��
ŭ=q�?��������?�Jؽhl�>�ݘ>l��#�@>gB�?L|�����ę,?���d9�>A��>���E`>���?R���|z��"Y?m���>�%�>�� ��f�=�7�?B/��@���RH#?m���U>O��>���'tP>o�?*����x��+?#*�8o�>X�>^�����N=�?������"?�˽�I�>�Q�>R��&�>��?���\9��Z(?p��2��>Gw�>���_�=�*�?>����#����?�!���2�>S��>����0>+��?��������C?3뻈?�>��>4h����=႓?�6���h�?0-Y�N�:������V��ݨ>������>� d@���?`w7�AM����U�=��>�,�=W��>��c@͏�?�"F��������5���>[�=g��>��_@M܆?�1��[��mG�!�=�m�>M1��9��>n�a@���?��:�N�����I�lO���>��c�g�k>f@�Q�?�<����{xE�җ�<���>}�=sI�>f3^@��?x�?�|�0��Z��u+%�;��>���<��>D�`@��v?Bo<���*��eὑm�=��>g�s=�`>�4b@�$�?�1����|n����>8K�=Aޯ>؆c@]^�?lF�n˽�7�Ҍ=��>=*Q=籍>��f@��y?�I[���м�ѽ��!=���>�6�=���>�d]@�V�?nUP���2�ɱ����}��>�#��+�>f@�t?"mX�U8*������z����>�I���bX>^!a@�v?��?��K@��9��&��G8�>��A�!�>�q`@2 u?HY�y���N�õB=k��>�&:{֮>?c@�t?�V�����|���z=��>�W=�1v>��^@�?_`����O>*����>�	�����H0>�q����>�I���J>N��7�>�l���1�d�C>w��!?&ѽ�@�>\�����>�ɾ��)�C�g>��r�!��>����22>�n�
�>g���g+�6>ظr�
�?_�%�>���F��>rоf���ae>�(w���>l��i!Y>��Ҿ��>����'v���P>Zkw��]?{�R��ep>���,�>S����U#��kC>n�x���??7#��U>ޭ�޲�>������8>��u�{+�>�)U��
�>$�׾���>�O�������>0w���?).��*�>���^��>�[����*����=�_s�`��>�6\�U=>�߾Ɵ�>�ξ�+�=��=6y���?��=�O��>����&�>��~����>|lp��?rK2��n>�2��4�>���q3�~�E>�z���?r���_>@�پH��>����1��w">*;z��:�>8�0���> {ϾL��>��;�}0�TO->�gz�\�?݈��k>�y��{�>C������>��x�UD��m�<*o+��B�GU����s����?�9`?�J���-=��
������76��/��rB=�\�?K�S?�L����=�����z�[�T�XJ����<#�?8Q?�L�8�	>t�(������O������H<"@�?��]?�fK�s%L=���@�w�-�m��V��H͊�?��V?&C���=$&��8��l�ڽ�̆�Z�|�?"d?L�A��=��!���M�wu�ރj��)�=W��?�pT?(`K�n>��������p��K��r78���?�e?�AK�QN�=m#��r�h��N_��Ht}=+��?�$f?P�G�aN=���}\��}��
w�x9c����?�kM?�=I���= �(��ǣ�B���JCn��b=1��?]�d?eE���>�c�9����D9��y��>�%�?9�T?p�E�#��=rh�Cբ��,������2����"�?�mI?��E� ��=.R�������������9\;���?��f?Z�I���=�<+���f��sX�8s���񜽚��?�B\?�L�W�=V�����?y��a���C��"�?�%R?jk1?ٍ�?��}?��a=�˾ۙ?�*1>�?"04?j	!?K��?���?
�=L���'�?�~�=<n?��B?Ծ)?c�?B}|?�A�=ͨ���?gPH=3�>�_2?F??W��?�!�?Y��=d���у?�GR>C�>l5?r�?;'�?��?�i�=�T����>�)�=���>d<6?�T?G+�?�j�?�l�<v�����>�H>�J�>��Q?�Q6?��?U��?��=$k���6�>|�>M ?
�S?�n8?��?y��?�'w=&���6y?���=f��>>�V?\�(?���?R΁?������#��>>��=Q+�>�q<?��3?�V�?-?��S��>~�3� ?�?>yi�>F7P?@w/?Ӌ�?Qf{?s������?���=�@�>.bY?Z-?�#�?WJ�?��L��V��W�?HE>W��> �P?<�(?K��?"4x?���<�O��v?=�H>���>��E?�|*?,��?�}?�E�@½����>f��=�B�>BGK?$v$?��?�߆?��e=�p�� ?&uV>���>>�W?T�6?���?���?u�T=�[����>���=1��>;D?�L2=�H>�]��%�v��ײ>�?���`@#y~>��=# >8]p������>5��?�����^@-��>��%> ��=`c��ꏾt�>Y�?-�a��(e@I��>� >=es>����uמ��^�>Ӊ�?�B��C�`@���>�k<��T>'�ad�����>�t�?qqv��'e@���>��>�bm>0��i˾pά>+*�?#����f@55�>�
=�S>��������t�>�;�?`����]@s�>L�>m>4����}�����>��?[���]@0hC>���=N��=J�c�ӡ���%�>�5�?�����d@��@>}�=�u>��C�&���ҡ>��?�p�gv_@���>��
=y	x>��&������>k��?��c���`@xu>��=�q�=����1>��̈�>3p�?C�m��Ec@��>]��=��%>2/��!�����>Mh�? ^�A�\@i�>@�<V@>��'�V��I��>s2�?�\���e@�[�>`�*>��l>�@!�b�|�X��>_��?����W%^@=��>��=��>�䇾S�ƾ���>��?@ʵ��e@�{�>$!,��������?@6$����?"ş?�(�>e�Ӿ�4�>��V��.�Aօ?t��?��?֣�?��>���T�>&:��v4�I��?L�'�?���?J1�>�wƾ���>?��]؀�it�?��$����?T��?R	�>)F�?9�>�YX� 6_�Ӎ�?#�
���?t�?�#�>M]ﾻݿ>d���vd��_Y�?�*+��ߔ?.w�?Խ>5�Ҿ���>�&�܆(���?ul�ų�?���?&~�>ߢ�W��>����m����?��K��?���?½�>۾���>�������?M��� �?�v�?Zȡ>%;�s�>6���:�P���?w �y�?D�?�Ʈ>�۾�=�>�b���J��΄?���?,�?L�>����C�>v 3�"`,���?�"��4�?���?���>�cӾ�R�>��jU��3�?���m��?>�?>A�>_�߾'��>�yv�ނQ��?" !��0�?��?�[�>������>� q���H�S��?K�m�?ޫ�?���>[��U{�>i���H)����?������?H��?���>�����>�cݾ�p@Ԟ�=_웾�lZ��A=̐�=அ<�P�����m@�/>����N�MP4=B,3=5j�=��&������m@+� >Sҝ�PwS�۳=rL=d�8=V��v���q@0K>젾:9m���=�8��p�;����a����gp@)A�=�鞾��N�g�=��=魹=׽8G��cl@��=qO��@'W�Y�^==��^=䆭�R��,Ji@�i�=cg��J�[��ˈ<`ސ=Y��=�֒��d�n@I��=�j��Na�,�>�H=
cV=���B_���p@:؇<'XھnBa�\�,���=9�	>�V>�4���Jk@�%>�2㾚=g�����o'ڼq��<*~��2Q� �q@0��=���D�[��T�<;�<o��<��9�(n �~�p@"��<m����X��|>D� �҂*=�v4�V��F�n@ �==̾>%n��i6=�ļfer=Ak3��:�vo@��f<�k��B�e���u=�&9=Έ=����� @q@8_\=�A��`�`�*j�:V�=�O<'��F@��/m@m�;�����dS�_R�= n�=�b>��-�|�(�u�:�6>��.�>*�@@74�3��y�5�*IZ�A�z��ۑ���S��.	?
�A@�IL��X	�e;"���L�����Q��cd���"?
I@@v��Ń���8��1Z��N��'��S?Z�/?܋@@o�3�MQ�e�I���Q��F���+=g�e���?��B@Wu�k���J�z�V�<G)��L=�>�)�?6�>@�5���B��\'��R�@𜾞^��[�=�	3?�f:@�j��l���?���?�q|�J���M��h? );@�u0��
�˺&�zQ�H�]�.�
<�]���$?��?@Q󫽡�&��'�^
L��3���D=�wd�=!?F�<@���u6�G)���f�x�a��<����?��7�>�B@�7�A�	�1�+�2zg�x�������[�j��>��?@�F�{D���,�t[�v#�ؼT=+�@�տ?LP>@��!�am!���(���A�|���P#?��;T�K?�&>@M�3��U�y�3�p�C��b����ؼQ�V�#� ?*cD@1n���o
�c�<��h�����bL���QA��?"�B@�LQ�7M��6J�4�M���3?�j>�F*?th��Qf*?�}��V!���U� ?5�#?k�>%>?Jݚ�]�2?���k��sm���$?=&?��.>�H
?�X���1?�P��ٜ�>y��?��)?G�>yp?Z�6�-�A?Q� ����f�^�N�?��,?Q1(>)?����W$?��vA�����?�1D?��>�,?�靾�1?:J���ۘ���Ὀ�?MU6?�}n>Ø?T�E�I�5?���l���PHo��?1z4?vV$>�?y,�U�!?va��隿��,��;�>o�E?�Cb>w�&?x����|-?z���y����c�4�?a� ?���>A� ?����k+?�+�xݖ��?�*G?��D?��M>( ?d' �k�D?� �ܢ�B<��@�>�h,?u�W>O[,?*jK�{�/?�y���e���P��J?c[@?��K>�/)?X�I���=?3��꡿^�B@�>_^!?E=)>EJ&?�E��om&?�%�
������>��;?U�a>-?7w���*?�������L����?Y�4?��A>+� ?|fI���>?,��&ĕ���ս~�
?KEƽ�o�"9Խ���?K^?1n�9�?�vf������Z��Zt�U���t3�?'{?P��T�>Z�v��4�k�̽��^��*R�� @�.?�3<���>X�R��Of�q��~+j����E�?3�?>���?��d�Ȥ��Q��:R�j{��2@<7?���=���>V(i�9]��D`���\��8L��	�? s&?��=���>�W����U�	��k�'��m�@�?��f<LA�>�V���m�/��M�"	#���?�� ?+�O��W?*�a����΃��fa��ֽ���?��?�_꼬q
?4�f�"��[O�l�l��k ��(@L<?� f;�?�W���f�3��x�i��ʘ�^��?FL$?T�=z�?�R���<�x����o����@@�#?�=��?��p���D�$���<)p�pЂ�Y��?N?Z��T?h�f�lPf������S��H����?k9?�v����>�V�;)��Y���m���F����?��?�y�=���>�u��fH���ΛZ�G����?�/ ?�v����>��z�+�j�8��<��>��u>'g=���?S�.�}��>c�e������;B��>�NG>��=$��?)]-���>�������҉�=M?�F�>�1>���?���|r>�s.�����~=fZ�>�?>)�>��?���R�>W�"�������=E��>3�Z>�|�=1��?I���R�>�6�k}��i�=}8�>2��>��|=���?.����>I9�����<���>(5�>���<���?#����>s?-��轿p =�o�>��>20>�{�?��-���s>���˾�s�J=`�>?<> S�=�?�?�n����>O.7�[�����:=E�?[&�>vT>,c�?]$���>���)���qMp=�e?eٓ>�]�=��?��
�,j\>M(�E���?~c=� ?V�>?�A>���?�r����>/J.�孿��=j��>Ɯ>r��=��?�)��ԣ>?�&��3����	>8G�>b�>� �=g��?��$��a>[�(�u������<�g�>&��>��5>���?uz'�AR�>�!2��N���V=ZJ�>�f>��7=\^�?&��>�3��ﵿ:��tY������� ?<!�?��>���>F�z>i����=H��u�U�==x�>�6{?�u�>nJ�>"�>�w��#�X�a�>15y?,�`>��f>1>.�f�uQ�<�g�Kj=5��>���?��L>�W�>׻U>��{��������A��=Ӗ ?�,�?�')>;�m>J�j>L`��ν�`�&܍<Wx�>UՁ?�:>�)>إ�>.e�V��{���A<���>_7�?�-�=���><8�>�-o�R妽�y����=h(�>jS�?�6:>y<>��P>��i��I��g�w�H;�B?�?B�D>%�$>u>M>��l�!���v��
�=x��>�݆?7�>_g5>+l�>\�����	=WD
��`�=��>Uă?�eQ>�y>��|>F@���?=����	#=�y�>���?�~,>m�Q>�<Z>7	��"B��c�����=���>FƆ?��>���>#
l>�]�����G%�$�L:z3�>I>?_�>;�>��E>.#e��o�����n;�?9�?D�=>�2m>�e>��t�Qn��%�F�����>]�~?��z>�C�>x��>�@��_�ک�����W>�{�����>���>}��>3��@�e�pW���S޾T#�>&���>';�>�ۓ>��@��������ξ�X�>iF��p>�_�>)�>��@�^������T��>�N>��{6>袀>8�\>�ۂ@3`��K����;-r>~X���jL>�`y>/\>��@�ȱ�Yq���پd4Q>b�M�,Z�=��y>/��>ր@Mꍾ:����F�U�>@w����1>���>�E�>gq�@����:���K����>�@�sK>}i�>˅�>���@,�u�:*����Ⱦ���>�ʫ���
>���>z&d>YK�@w��|L��|�	��ہ>L�c��z>UΩ>�{�>i�@���b*��y���@>���3Pj>1ٝ>Ka�>[<�@s�����M�k �(��>4@���X>=�>��>��@%d��Z���(���2�>2`��5�>��>!r�>��@�o�L����,�X�9>�@O���;>_��>�ù>	�@a ��\��F׾ιv>�(��9��>K��>��i>!&�@ge���U�o�Ѿ4��>:���>��>�/V>���۾���?ȫ�=���!�Q@���=ğQ��R?d���޾�k�?��C>��ڽ1�M@�>U��?DQ ��
�O��?h�">t��o;S@,>0tQ��%?(Ͼt���U�?R�>e�2�۹O@���=)d��c%?����%˾�p�?�
�=��s�I@���=��?��?]ھ~��_O�?"�=�䷽1�Q@.�1>����
?���H�Ѿ)�?��=�?��&L@��=����<&?Zg��
�C)�?�S%>���&J@�"�=���g*?��ھN�����?�W>>.0���K@1�@>��=��$?0�־v�����?��>$ᑽu�S@E�=�5����	?�vƾ�3Ⱦ���?f�#>���3<P@ʇ=���A"?�bҾh�����?bL,>��$�݆P@z�D>��ý]#?hоZȾ��?�7 >�a���S@S�2>��>��y?�;ھ�x����?��>1R���O@��>fA�s�?�.پ~�ѾS��?�.X>W��7R@C�:=ۢ��I ?�U�|%	��F�?x-�=;����K@�53=X�A�9m?y����?8�d@.v�<�ὟB�&�O=�#ʾ�%�=��־Գ?<e@�b=�c���;��*�<��ž�4�=dUվB{?FKc@�M'�8�%�5A*��ZӼ�բ���=�Kƾ�?R�c@�������Ѧ�Z\�=j��q��<�Pʾ�"?�cf@	c��Z�&��,��|>ݾf->�l۾�T?��g@ۨ�=1�S�(���� �ƾ4��<|�о�D?��^@��!=f3��;&���=��� ^>t�Ѿq��>|=g@�!�;ȝ�AL(����<D����=b��;�>n�c@M�<LY*�q:9�`&=�_��\�>��龂?�f@C �;$t���&��!�=�3��V�;:���1�>�Gb@%F=�gٽ�[;�T�<�j��1N=@r�O��>��a@�7�<l�3�cV1�F� =��;��;=(�Ǿ�?X�c@M��� P�'��F��p���R��b`���t?p�a@۸o<��&�#�H1=аپKg�=�����?N^@���&�E�ߢ5�)��=�þ%�=�'�l0?d�`@�d=�E��[M0�΃��!d�=	@��v?8*>��S[?��=�Tٿ����	iL������?�h>_���rO?�B"���ڿMp[��@@�G��)*?Da>3��hO?fÂ=#9ܿ�����+J��࠿��?ז�=A���C?�'
>��䉴�iE2������?a&|>0�%��k?wf>7��������1����oN?��=h�
��k?ڛ�=�6ٿ�㋾ekL����B?�k>���9C?Y|�<Ǖ�(H��af<��u���?eb>*�#���J?��<�n�l_��_�)��$��� ?��0>���ork?;H>=���̤`��*���e�?�%O>�6��SM?��=Q-����H�E���/?E&&>����`?ė�=�ӿJ�w�K7-�3y����?��^>����)d?�l=i�ؿd���߭-����I� ?k�>(W%�k�a?�� >C�׿h˛�9�0�+ɟ���?��Q>"U ���M?�J=W�ֿ<�SE%�SR���?��F>>8&���c?����Կ �m���(��v��o�*?��6>9���H?��>_<�m8m�n&���'���/�}I����>۹>ŵv?ð.����>���?o�%�>S1�N);�W��>gD�>��?��,��6 ?�N@o(���ۂʽ��>7U�>ڔ�?�9�_?P�@5f+�׆��ݽ���>��>�E�?��B���>�~@7a#��&���ӽ��>��>Te�?{�@�Cr�>�6
@-���6.�;�w�>��{>�֋?C�I�/��>@2
@���^�*�}��T�>C �>NV�?_�=���>@�p��6�?s�����>?�>!>�?�B�XT�>b�@=-#���-���Ͻ7>�>{S�>�r�?��M�r��>n�@��'�2T5����ë�>��>j��?QcB����>d�@�;+��n�9Q��G�>c��>c�w?[LH�~�>�@�Y �K]���9�>�V�>�}�?�<��V�>�� @�2��1�~�)�Ǵ>�>\w?5�.��=?��@'@�
16��?�ן�>�T�>��?�+��'�>N	@��#�r�6�-yY��B�>	>�>�x?;�4����>D�@��0�,0�rR;�	�>/�>��?��;�gA�>MJ @��@��w?.�����U�����>:>|�>T�A���"@˃e?�!�1�"�����JM޾�H>iE�=��O���%@�,`?ٻ���(�k.��%���9�=H>�<��P� i!@��|?���7*��ޱ�����n�5>���=�B:�\v @J �?��:�ߜ&�`YH�V��9�#=l�D>�YN�|�$@{�w?i�5��������w����C=&�B>V*,��R @��z?�2��Q"�qⅾZ��x(=4�?=�U��.@�O]?�7��=+��$g��侕D�=�~T=$,F� @5~e?�8�qs�矑�v/
��=��E=n7�6A@��u?��5����!W��]���mJ>wD�=֚G���!@?�Y?�Q�u��g钾�;j;>���=
P���@{zW?/��A��m���ui�3d�=A��=�}F�ڌ#@S"t?ݟ:�52�2�v�h�����=�=DI-�>@@�?Y?�<#�eR�F�������>�U>h_I��@M_?!��_��D��]����>�=(>�;A���%@��?�."�UE��-o�S�۾E>Y�=*�>�gI�l��>Y<��ޢ?y)�=&*>�G� 3�?mY>S����6�>����f�?��2=��>Wpw�?��P>[Ժ�x�>�r��Mk�?yn�=Z�>��Dܨ?��:>'A����>�^�!�?���=�>���|ܬ?�q>��7�.��>����7�?�7>�/>e���?��>f*���b�>4v�Ю?(��<r>ɑ��T�?� T> Z����>�����?�j�=�I{>y�˟?/L�>�b�hr�>����M��?-�=̩x>�������?��s>�½�>+%�1g�?�<�=�]n>ә迸�?�A>qN���>q���ݢ?�0B�6�>���6��?��>Y�.��>K��ء?�bp=�k>���?��*>����[�>)��K+�?k��=A�U>�1���U�??�>�7��&�>>3�!ѥ?���=8��=�%�؉�?d�V>c�J�P<�>������?�c�=�C>������?��>���K�>O�6�??+�=s�l>�J��po�?t�>���p�>�1��m�?�U=a�+>YJ�����?�J0>��=(˾'@��=^��]�>�>;@^�Y�?N_;>�����@��E>$V���?��=�~�F�?�S@>l6��/@�{�>�>
���?�1>/����?&�><cվ�@���=n�	�JW?�=����:?y��=�]���@i�b>���4/?�(>�?���>�z@>貕�e0@�e>�����?��=��͌?J�=By��I�@��>�7&� H?YT>��C��?!�=J�˾��@�yQ>�!�t?�@0>53k��?-x�=�ʖ��;@�U>0.�GK�>��<>sFM��?c�=�[����@�0M>����v?+��=i�y�C*?4�>>�'����@��Y>�O*��
?妚=�/)�X*�>�j>�����b@=�X>j8�7��>'L�=���P ?}�=d�ؾ�@�k>fV	�T�?;��=��z��?�4>�׾U@cls>��"�x�>��N=��L���?�6�= ���+.@Qtx>�,���?�i=s>�C�?EM�=��ž}�@�>�J(�� �>�6">aK��<?��?0�?��@i����/��->{'+>�HW>2�>=M�?��?��@��V.�ɜ>�f>�q=��>��?�e�?�u@�N��1U"=.�= ��>Xlc=fT�>� �?D��?=X�? ���n���Ï=r��>�J>�Z�>���?b��?Zm�?Fl����=w�>>�>&q�=���>���?�Ǥ?�*@B�a�UO��
��=M�>��>L��>a �?���?q��?����9�Q=Z��="\�>�}= x�>�r�?l�?��@�{_��7�<<
>QQ>��U>5�>���?��?�@�a��A6j��</�{>�K�=|��>�w�?�
�?� @bNq�N�n����=��> >>�j�>�R�?���?@�f�Am<>��=�>R=9>�:�>�(�?���?��@%��#0<�ք=��>IS�=��>o��?���?/.@D��B�<� >�n�>e�=���>���?�җ?�)@V�>��U��4�>��E>^u�=�~�>���?b��?o��?�З�˗/=�ܮ<�[>,$�=��>���?FҤ?ͥ@�R�!�[�Pe�=�a�>/�=R��>/�B�&�>)���Q��N�n��9C@��ž>_�=74"��<$��@�>u���D�z����K@��ľt��=�&k�=�A��{�>t.������0C@\�ľSƈ=�{���7��&�>�(*�O��ǽT.F@�������=����kZ�O�>���.�Rs��l�D@�0ܾ�>�=�ƽ��w�M��>������>�ΑE@����r�UjD��t����>�������H�.�,�E@T|����=��������>Ԫ�b��8����I@�>��:�=����|����>��v���!��jἪ@K@���[7�=g�� &�Kw�>N칽UN��;�`B@�7�e�=��Ľ#%�'�>ěd���	�H���D,B@�X����9=��b���o�1�>&"-�	}��:�9t�G@Ĝ��>�A�����Û�>����R��;��#H@`�����=p��K����L�>��I��.��/޽>J@��¾Z�=�TQ�������> ~T�=-	�"�	���B@|B̾��7= w�3ކ�UH�>rQ�q�%�ҋ)�N�K@������<ǫ2��w8���?�-?f2��4���Hw>0���I@��K�"m���[?�~3?g���Ŧ�bt>h<ʾ
@7�]��T[��n#?��G?�������$u>@��8�@өP��-���?MU;?��L)���o>�����@!�?��X���??�6?�)�r����>�ɾ�`@�IY�/���[?��-?#�!�hҜ�:�}>����
�@��A�E	�ך+?��A?�'������=!A~��n@�JO��}@���"?�)4?��1��{z{>���0�
@S+F�y��1?s�.?Ű!���Y�K>D䓾��@�\]����%P	?I�A?m�����!j>�Ǿ�@�/Z�k�q�+�?s�0?}�+�B����]>�W��R�
@y�R�eN���?��5?���ݟ��>+þ@�Z���D��f*?G�F?/������e�"> R���y	@�WG��6�c"?�s)?k��B�����>4����-@OP��^m��2?�r4?���V���q�=�<@oaC���O�mW,?��/?�*�����-�=ސľ�@-�G�NM�>��ؽ�>=���>��=��L=v����d@:? �>��?����M�>�K�=��&<R��ʊe@�C?0?�>$9��y�1?���<����%��hb@b�?�T�>�a<�H-�F3?3�<P�;=�����c@*J?Ќ�>|��7M=�� ?}h��I�=����8�g@��?JT�>���<�GܽwR�>��<�������c@�=�>���>Sq?�(������>��b=4D=G�
��?^@�"?�Sw>p8��SI���N�>��<t�=�O���d@�?D��>�Y�:l��)�>�0�=+5ּi��p�d@�/?�>�o���H=���>�H�=a���g@�?��>]5���9���?b��=�5*��P���g@�,#?X%�>*�j�o�L=���>�(=�xo=��߾�^@��?��>�V���o;<"��>��=���<�/����c@� ?my>�ٽ��=�K�>���=-��=8ݾ�f@��?2%�>t]� �ѽ���>,=�[*�����`@��?���>|:˽~�н>��>��H=�Y����x_@�#?"�<?lPW>�Ⱦ{���gB������-�?r��?i=�? 2?ت)>p'��J��?&F��j�����?��?���?�O$?���=���=2��^�����fѢ?�u�?��?<z3?8>Sw�yL�I���׾� �?pF�?�$�?V�6?=�>�~ھ��"��9h���Ծީ�?�^�?���?�&.?�^>�����7�S I��\¾"n�?�M�?�ݩ?�d.?�8�>]	�%0Q��6e�aV˾x�? �?b��?��3?]�}>���l�G	B�I��BQ�?vަ?o��?�� ?�t>�{Ҿ�	.�yOS��ʾ�@�?�<�?��?^�8?{Շ>(��G&�yBR�aɲ��͙?:�?���?��H?�>�>~�Ⱦ��>��X������?"�?�ޮ?t�6?9E�>�		�M���H�?s̾��?"?�?]��?��D??A>�E�!|��})I�I������?��?��?̕5?�>O>�ھ��n�5�a�a+��?�ƚ?��?�tB?L�,>`ľ}*����[��񩾾�?Nl�?�U�?\^<?Ȕ0>zZ�K�/��d�G�xܕ?v`�?:��?1Iþ*�p�����Ep>��'?�[�?}þ�p���(�=;ץ���K��D���%�=E**?�,�?�~Ҿ�鰿���=��˾O"����˾���=�?��?Wo˾L��� �=�����o��A\ӾoMa>\� ?���?mξ2���a�>񚰾�,�ץھ{�>K�?��?,���d��?�=��Ҿ��{2˾sy>S�'?��?�뾐9����>�'��N*�����X>��?���?����'��j	>9e������V���">�g?���?�{��P���,>W���t���ξ@>e?�I�?3h�n�����k=��پx"���p��ȱl>O=?S@�?K�ʾ\���-��=U[�(+^���ƾd
2>!@'?�?�_Ͼh^����9=���VJ�K嚾V�R>�
?�2�?�;�������=+����b?�}���Q�J>�?���?)�Ҿx�¿��8=����(������ >�E?��?����qſ�+=�1��Z����ꩾ��>�?��?g��T��!��=[��V
N�i[���>�+'?3�?X��k����;>�X��f�??߿Tÿ�.{>�x?Ȃ�G��"��>bB��(@Y?���._�� �>���>�Xy��뾖"?M��h?�r���ʿ�#�>��?:��a鰾��>����Xi?��忂Dѿ��>,,?D,_��>Ѿ�?BW���lL?&鿔�ſ)�>���> ���J
?�/1��g?�����˿?`�>�o	?2�'�ƾ6Y?�ף�btR?_�迲�ſ�l�>��?갽ɦ޾�� ?Uu�HA?ߞݿ�6���.�>�`?�
a��bھ���>�D��N?�#⿤Ϳ;��>j@?Φƽ�����?xa����b?�V迤ȿP>�	?8&�	¾�q?Tf����E?��ֿ,Bȿ���>�%?����O޾n��>�*��S?�v׿g��[^>H_$?�KN��d����?$��;F?aIٿ
7Ŀ7�f>$?��P�2Z�����>���h�T?͎�VY¿���>�_?�GR���Ͼ
{�>U�K�4<\? ���ɿIEQ>��?p�8�>��,�?&l ��f?%�TпU^�>��	?�Lm��ž3R?�
���o�>�KL=��L=�������G�	$����#��t��?>k`��࿰�J�0��������ί$���(���k>'�̼AP��Ӧ]��lѾ�޿���X�$��o��թB>�/����<¥�le�%Y�_݈�X�����KG>[Ek�L�����W�����ݿF0����&���+���&>~�1��#������	�-9⿐ф��r%�9�z�{-[>$Oh��3w=$8T�h$Ͼ%��f�p�$�,m���9R>/ ��g��?O��oҾ��Q��Dg$�܁��Ty�>��_�j��c;��wɾA2忏���Nm!������/>ڟ%�����y���������e�f�'��oG��r9>��$���%���;8^Ͼ9�ῥ}u��5 ��0��Ƙ�>�O=���<,A���Ǿ��c���!��DV��Z>ˣ��ldM=�u�;�ľ-�����r�"�brt��NP>��%<�w�������]�߿����}(�����<J>m���b��<$��/ƾ=�����&��8���>����SD�=W� �Z5��L�m4r� V(�x2���T=�>��>�?]���?�MB�>��h��=9b�<��=؄]>�$?�6���'?_3B��c����<�ș=>�=`�G>_�?��Ƚ|�<?�D��)��P��ԉ<�;I=x�F>�F$?N�ὢI4?��>��e+�7���8��*F>P�:>�#?k"R��X<?�7E�<.���1=Дe�_��=��;>	�??� r3?�F@�gf.�<��<�2��Q�%>�!�>��?D���6?WE����4V�=/��N?>���>��?�3j�f?��A�#g&���A����*�p=l�>��,?m�ҽH??k�F��]D=��7=)�>�a�>CI ?:B�>�?_�D��w&�e�̼S;�=6>6��>Ǎ?���ƴ:?��<��$*��T�<�m"��\[=��>m#?�Nҽ��1?�DG��U&���=��Ӽ	ҷ=�,F>��:?D%A���&?knB�g!��5.���
��>�>>�;,?��6���%?�@������r�-O�=)b�=�ύ>��2?�\��X5?��@���%��e�л�,>���>�0?�Aٽ��6?�F�9�#��>���>i3��>�>�AV?#om��SU?�@��'?=�>��>�K�<_��>��k?-��4??O!@A>(?_�>�K�>�����>G\?�d��ER?�'@��?>��>� �6>9m?�8��N%C?��@yT'?w'�>=ձ>�n���]>��q?�:��қL?w|@�/4?}՜>c&�>Jw��4>G�d?a���7S?�C@��0?f�>�4�>�R��t>C�\?"}�xrL?�[@�t3?���>UXw>@�h*8>��S?@�N���K?e|@��=?�U�>	Š>����5�>� ^?�嚾�-H?��@�31?�*�>K;r>`���x>qcd?
�f��0K?�@ya<?�K�>�!�>8L�<>�ll?1����[?%�@��B?S%�>;�>�2����y>�;[?q��� cW?�Q@��:?1X�>-�>k��<�Ui>�UX?9rI�*�Z?��@	x+?���>��S>�Z�0�\>��a?���l�F?�K@w�?�>�v�>����Ӕ>![m?8�_� �G?ǃ@��-?%��>�M�>�������>-`?	_V� wB?�V@�%A?�-�?�<��u��<>U�>PΠ�%::����?W?�>n�D?3�?�z�=��=���>�s)��" ����?=Z�>�21?���?���=n>�k�?z^�%�!�sE�?���>�=S?7K�?���t��=��?���m�"��&�?�*�>�2?AA�?F|=ʡA�!�?��\��,4�m��?w<�>�iF?I��?9<���=$��>�'��ͺ3�Kr�?9B�>�T?�K�?����=b=ё?�p��#&���?r��>��Q?K�?� �<?���H��>Py˽'.�5��?[�>��M?��?��@����<EF	?:�B�߷8�k��?�E�>v7E?W�?��=�ә=�@?����i7����?[Q�><9?K�?_ޏ��p=�m	?0E����4�M�?�;�>�KB?'��?��ȶ��?�ȿ��,��c�?ӝ�>v�S?�?he=��=�?��=�Q�*�C��?�C�>�&H?�+�?!�)��<��?��|�ǫ5�?�?!��>n�O?��?��=Oy�=v��>^(Ͻų�i��?�,�>4'+?�m�?y��;r�:���> ��j,��?��>,�,?�ʆ>�w��8�p���ʽ
�\��;��>��q���A@7�K>#w�D�{���Խ�\��I��h�<a�~�S�;@��g>)JZ�Su������^�U1�a!>�$w�	o@@���>[C+��>��N)����S�R,��F>S�g���8@��N>��Q��r�����.:�����j�=63��7�?@>Jٙ����� �<:A�,$��10�=�u�@@#�D>�!���{���νސ9�
_Y���=�h��^=@�Z�>���x3�Z�Y�ؕZ�K��u/=�n��n>@�>�_~��TI�*�
�E��C<����=ňv��LB@%�:>Ȭ����/�3G�H�=�o>����=�}n��]>@e��>Ɉ���	-
���:�~KQ�E��=�|�5:@"o>e�C���ɗ���_���t�E�=��f��@@㝠>q�?���D�BS@�p�A�A�5��3�=�Po�U�?@�8w>��G�T\:�y*�r�D�@�>�Q�>����=;@=�7>\�����Խ��O��_߽lJ=I(g���9@�OK>�O�o��)��8�:���C�8�>�l�W�A@��7>� �>e>�?>��\#��HE��a�ޗ�$��>���>h���	��>��<�v����K���j�|�����'>�j_>���e�>�~=������Q��Ye��ˍ����>�ő>�(=��>�� �����-�Q���c�,���Z(>��>Ȯ�=[��>��W�����{�l�
yk�,������>T#�>���=ޗ�>��
�%���V{���ta�< ��6��>�XV>�C�=���>R�<����;���N�a��<���W�>D�>��<��>rY��)ݾ��S�p*d�<�q��p><��>�򑼗�>�v������&�"i�
Q��<�>��>���=���>wƕ��>��y���D�i�����/�>&:�>��R=���>�N�;��Ǿ�^�~�j�$⳾\�*>�
^>l��=}�>���0e���Q�""k�0���x�A>hf�>|�<���>yN�뤾��6�7b������xX>,Ƥ>*�=���>���L׾׿b���g�ľbDC>��><A=s2?�������!g��캾6_�>�p`>��=-��>�}�;݈߾+䙾v)k��k��yc?ì�>��>j��祋��J��CN��l�=~ƣ��5u?��>ݔ�>�v齷��wZ���̼	�>�H��o�l?��>���>���ҋ��RQ�13�]�>�D�`؃?$$�>ː�>�@��s��{V�TԾ��L=9M�� ~?̂�>;ͩ>%*�#���<L�������=͡��`hx?>��>���>�8�CO����\��'�?�g=�̾%r?���>�"�>ԕ�� ���c���Z��1>�ž��q?
�>w��>�Di����3^�u�|�+>�P۾�Tx?�A�>KM�>�q������0C��
�=m>����<g?�y�>'ñ>^�x�yr��+�N�p;���E�=w��OHi?$h�>cǾ>M�o�����EI�ƶ�4��=���@n�?���>�&�>��m�k���=HR�ku���>w����h?��>�
�>
��Ӌ�+�\�"�߽"6>ԡ��&e?��>� �>N6��,���bT�QN���FQ=a�ܾ`?��>�}�>��S�K���?X=�UH	�U*=0���#l?���>��> q"�����>V�Z��K;>E�g �=�['>�|˾h����3�D�.?��>#-O@q�=)T�=-3e>v��*���Ǒ?���%?c��=��H@`�'=�x>%�>��پ�qg��/��9&?� �=�PI@|8>�c->��5>҈վ�a���,���?�
K=��N@;$i=ew]>c�=�������4�H$?b�=i�Q@�'5>�5>��m>Fm��š%�748��H?�ø=��O@��2>iZZ>'<>l6���5���%�HO+?*>QQ@�a=M([>��D>��ܾ��-��+!�J�+?(�>-�Q@��=M-*>�q�=�����;�Ӝ9��$)?��+>u�O@z!>��S>ϖB>�۾�5�=q@���?$�>�`I@���=�S�=e� >���]�#�!M7��.#?��[=�I@wY=�lV>�L>�۾i�/���)�x ?5>eQ@���=g�G>[��=�;ƾq�&���:��m(?�~>K�Q@a�=]c>-�8>jmȾr���e ���?>��=oJ@H�I=M�=��=>�;��V�kp&��u*?OK2>P@\�{=�2>W�">Ͼ;4��8���?��
>	�I@�^�=�&ľC����$�o@?�V��KF��iy��G@���<9T��*�@.�cy?b`۾,;���Ǉ�e@d�=��ʾ�r�m7&��?�L���cR�����O@$`�=���z�Cz)�� !?2Bپ�2j�rr��6@�R<	���S���)���?�����{��q�O@��)>�Ӿ�޽U�&��?����z����m��l@�>P�����1;)�5?t����	v�v���	@6\�=j���;gY�6)��?�����g��q���Z@a�>?H���f�H/�g_?|ӻ���6��7��_
@�o	>�0��O�B����۳?0�������W�n��z@�`�=�A��gy1�|��y?:�Ǿ歌�0т�s�@X�w=������ ��'#?��վ�~�����3r@��=Q�ȾC����"���?��ݾ亐� ���+7@�߸={{þ��h��8"�W�?6ϔ������~r�/n@�)�=��"��,��Z ?>������v�3�@���=�#¾�?��"���?Ɔ���d��(t�k4@��'=���>j�Y��gw?�2���⾛�(@���>=sv=��?¿�>�S�댅?�t��Ծ�0@�>\u�=���?}�>��V����?M���N��A�0@~��>�<M�?P��>
�R��S�?�>��Z`޾�/@���>���=+��?z��>�F����?dJ�x���5Q0@�W�>�A3>�1�?B4�>d=�)q|?ym��LΕ��2@x9�>�l>e��?DB�>�-;��ĉ?�BX�T����x0@x��>��=M-�?���>�N�`L�?)K�����'m.@H�>M�=�y�?�s�>��D���z?�0���k���%0@��>��=-��?2!�> bG�(��?-����þ.@.�>e0>�$�?2đ>��a�i�?�|������|)@&��>�>�?�s�>x�;����?G嚾�d����-@�-�>��=��?R�>FT��n�?K\��r׾��*@���>M:@=Ww�?d�>xU:��?j�C�:GϾ�#-@�!�>���='��?���>E��2�?��X�殾�,@���>Η=m~�?���>�M��+�?p������`)@L�>IG�=٦�?�)���g=�q�?��Z>�C�<4��=�>�9��<�Z�>��5�6OJ�i�?y<P>��=f�;��>�h�<�>9�,�I�ν���?�$>�e;�.�=��8��a�<��>�]7��ɽ���?y}(>�W��;-�=ܥ<�.RT=���>�,<��
����?K|�>�u����<'>�T#λ�9�><������ٌ?��>�#:����L<�m�=x9�>�,��%ؼݮ�?a�>p�=���=��8��؃=P��>)8��'�<�/�?y�S>�(�ڳ�=^J8��=�>W�+�� ܼ��?��>>V?V=���=t�@����:U�>�C��4n<5l�?UT>��_=�Q;�E��剥>#�.�ʣ<���?՚V>})i=�<�<&�9��ێ=z��>�?�t\<���?��>'�n:t��8T�8�!�!����>�n)�Fn���5�?̀>������=��>����Y�>g�#�A@~=��z?�f8>peA�'
�n�7��}�a��>�#"�k�#��?��>.��*��< �<��;==���>�0��Ы<�{�?Ӷ>�9�����-<��;H��(�>��>^�<���>�����p�=��	?����@�O����M%>�=>��>�N���>(>w�?�h�
,�	���L>Rs~�-�R>�R��	�>/� ?~v��J�A1����S>��K��U�>JO�Z�=��>(�p/.��W�$$�>�30�?q">�o���r=l��>5`�=y�ix�m�>0�
��>�����=��>�� �QG+�����U>xc^=��y>�e��}q�=���>T���-%�!��o^3>����(*�>�
 �!�>y�?�����-�ߥ���2>��<��>��=Ê=��?��n[����_\:>^�<��>4�=025=��>,%��(	�=��I�>dm��s�'>R��=�*�=��>����3
�σ�ȕ�>=��;d��>�/����=ܛ�>ce��+ ��C�����>H�M(3>)����p=؇?�$ ���&��h���>fb��4>���<M�>̳�>:��{����6[�>*h=�?>񻹼#�>R	�>�r���!��g��	�>����I��> ۴=C�<��>B~��x�k���=�>m��j{�=�X�����>w�M��)+>s6x�Hrs���k>D�j����=V�P�?>F�҈)>��H�v�w�KF�>C'ǽ^4���ľ���>)�M�
Ys>��.�	i��^Q�>���b�&=�*־��>��M��>����9��R�>;��a��ɾ�#�>�oN��8!>9�S�E{��1�>�˽{��=����1�>��O�2"1>0�&�{�A��>Q�Z�{I�=>�׾��>��N��XQ>�����F�f>�՜���#=;���) ?�6L���%>w�_�1ׅ�/�>I���'{=t��r?UhJ�h p>	���뮍�SC�>l1�	�=׾�:�>�2K��b[>�%�w���c�>w�:�׼�`����>LM�� >�)�{���(�o>�7�����@k�����>e,K�X�#>Y�G�q�y��ٙ>�?����=��\M?�(M�'	>�	j��}w�34�>�)<�hq6<��ʾCk�>u}L�a�>�8�Ѕ��y�>�z��`�κ2����>�pF��'>�e��e���k>P���K=@>����?�N�� �>��g�J��S/�AО�-5�i2�U�35���ս?&�:8S*�G�.�̠���������!É�HgA���+�Sb�=nI�O�N�{����m�������
cF�%�#�d@V�d�C�YBH�������(��;��TnQ�C�$�Y��;b�>�%9.�y���)i�ˏ�����SP���H�=N�*��4/�%����|���j�G�+FK�Q��=�A#�5�3����yA���P����v�,�#���a=�,'���B�]�����:��Rn�>�.�OW�ƛq=D/6���B��h��Kg ��d�턞��H�1k�����(2���/�̜��s�u+�[1��*�-��U���Q=�v@�o�?��������� �����B07�s��-��=��$���O��m��6l��4�����;A��ǂ���=��;�E�T��`�������Q�������7�u���\�&���;�Aʞ�:'��]��̵���;������=�O7��P��n����������*)4�,}�^x@�j�C�#lR�u���.��3��	]����/��꺽X�>=�/=��NA�?��:PLp>4+�D��&E�> ����%>���<&��9>�
�>~ -�Uh�*3�> ?��,jv>0l=1=��K<��>|�0��j¾�J�> ����Q>�-���A��B%�B�>�*��Ǿ>ۡ>F���P�=�C�=�y:��x�=�C�>2*��:оh�>����� E>�#=�:�GH�=�g�>��.����t�>�A��pc�=��S=�m2�4�>��>0�0�ؖ�2��>�&��NYz>.�=�zE���<�8s>,)������>��tV_>����oB�� 9=N�y>�0��|񾰼�>�'���-�=�&�=�Z'�_�N�%�>��0�mʾ���>�J���e�= �:��8��
�=�z�>�,/�_����>4&��=��=M�F��:�H�o>��-���ʾ���><Ŧ� z.>�jf=UK���=��>d�)�����:�>T秿J�`>	S �W�I��-�
�f>��-��o����>T*��إm>b6�i..�̹>ʇ�>�E-�C¾DI�>X���6�>���[�$���>r��>�C,�����>�E���#[>7r;����YZ��U4�8H���Z���J��
�n�|K��i��y��\s-�x)�w�y��#?��>�e�.�ϯ�%��M3}�*[���X��;����S�.���㾓�����x��r�ȓ��Mt�>�C�����z,����Ƙ��7����#��]���]�65K��&�q5/�my��w��r��`�#�� ���u��IM��5�7�0�������+ې���(������S�jA��-������s���Q���H�$����q�m���O�	����)�r��'ľA�z�l�(��O
�9Qd��J�VB���q���
�����rl+��c����f���U�@��h���������E萿Ʀ7������m�$�;�o��1��`�������?���3�*��-a�<BD��
����^f��[���a!���7��=��5�y���Q��C�]�2�x�������x��x �a���Ic���5���������
�����9Ay��2������j��EB����}b&��L���ξ�ǉ�L�(� X	��fr��E@��[�������d%>��>��"��?XW\�9��>���?���2�?��&>�Ew>�:���c?~�V�m��>�:h?��<	�>r�R>i{0>�:�gS�>�y[�9��>��j?x-��)�?[��=�� >|T;���
?�u[�}��>`�?8��ă?�с>�Cp>��@��?��^����>8X�??�$�?\�	>�:>Z<�?й^���>�Mv?lh<�!?��2>��S>#F��?�[�%��>_Kx?*ޙ�-N�>�Og>�>��<$�?�{Z���	?���?%�l�?���=�P'>�<��,�?]��:�>��~?���*�?ӟ>��^>�t=�>�>�]����>@�o?��ռ 6?�M>���>m��f�?��^���>�7�?�)����?�O2>�@/>`����4"?�W�-{?8��?m�M���?`�>�x>�b��N�>��X��`�>7w?4ސ�ϧ�>i�>�eL>^i{� ]?�X��y�>k�v?�!ϼJh?L`5>� q>'^��h?�>`�å�>�r?��Ƚ�q?׆>��	>�Os���?>&\�+q�>rxk?�56����>��L?_����s���a�����Z�!>6�!@0�f?Ɖ?l�??!��]���\'�Hj��^I=�� @ D~?���>8�F?+፾,hl���#�������=^&@���?$ ?�gF?��̾����.���ws���h=��%@R\s?���>�;M?Q���Є��}&��,�P��=Z�"@�z~?���>�	T?s�ھ����4m���께��=��"@2mr?�`?��9?��Ǿ�?��`�u��6ۻ@�=h�'@��o?���>|K8?U����ZB���[�F�ý��=@�!@8$y?���>�8,?eܾ�(V��X"��"�_i�=،!@�t?BD�>{N?����C���TM�����'�=ި(@��}?�o�>�70?ug����E��i��&��8�=�1(@g{?P^�>�5?G����X+L�T�Z�2��=��#@���?�5?�	,?�+��;z���h��tM�"˥=�f#@[�?���>�QP?;m��cń�1��D�����=��%@���?���>D�J?����Ί��o���Ȭ��|=L�&@���?a?^�A?���׬���6I��&;�1>r�!@.�a?��>�+�����ǎq�}<��aA��~:?&�?�>�b���#�Ͼ�#N�͊Q��@���0?d��ь�>�Ja��2�G˾���N<��C�QI?�=��QB�>f�3���=׾M'��wV�𽾽T�>?�O���>��a�~���ب��.���B6�qS:<��5?rǮ����>��a���]�A
���б�R���;9@@?*���{�>R�d����������+rJ�-`��V�)?r�<wV�>��`�E�2���������{Y��sd�gN>?������>�k`�+���y���p��I�H��o��>P?>0�s�>J�a���|��̾Q�P���O�����;O?�z����>L�b�����I���N�J�X�E�R<�)?�ﹽ��>�G`��70���۾�����4K�4�	�@&5?�����u�>"`���O�{Mоm[���bH���>;�7??�����O�>{^�-D@���ž〾)�H�7��^0?��b���>*\�D��i��r�c�w�L�����F3?�C�YL�> h\�y�G��>���G�;�+3<�oC?<�%��>��d����>I ?��?��!?��������=?�Ax��>��>;��>ӟ??��P�X� ��TT?��4��F>��>��>��?v]?��A�6Q��:?|���/#>Q�>I��>O\,?R��>��ս?��g^?%�|��у>��>E?�>�?�$?}�u����I?���X��>�
�>s[�>W1?��?YF)����g�D?�EH�5>uĘ>�5?�?��?J�J�A??pK��y >[��>�f�>o�#?��>�K�d���_?�EE�'�s>s�>}�>�+?�4
?��x�,� ��	_?����E] >գ�>1��>��1?Z?9K�r8���H?�bX�Ϯc>�~>���>��.?2�?���P��;L[?��[���d>q�>!��>}�?��
?� H������N?�?r��}	>�1�>���>��!?	"?���x����Z?D���Ղ>���>�D�>��?:^�>Dn��x��5iI?$L�x(>J�>�>�?�b?�R�:t��H?��h�b>-G�>�J�>N\	?t'?`:��<��q9?��{���>�;��Z��Zp>I���"x���S>Z@���߽)���N� �v��8�>�:��p}'���8>�<	��������S��坟�@''>qX���>H�$�i=7����/����=���ʒ���<>M⥿DdG����=�q�ڠi;$�0��. �Pnn�Ɛ�=;h��~_0���>��
�~ ���1�=�����K�ϑI>����=ҽ1�>4�������=d��8��fzX>û��q���&κ=������?I<F7��W�*��=������9�5>���{��� �={l ������N�=���$�r���9>���..��&/9=����Т�Zu6>�᱿�/)��>��������2=�D���"i� ��=S����B7���>�/��e���o=�����h����>�Ū�8�P���=�s��ƽd��=/��Hn�6�8>�ܮ�6���Qe=ғ��;ӻ	��<}���R�?��N=��������=�9��6a��|����y_� �>}B��dA ��S>���x�RC�=����HU��:D>C㱿ؼ�����=��	��v��Y��o�)�:�>c����2A@@�>���:6Ǝ���?Mb ���>������LU@@e�>�+���p��>�]9����>7 ��+S���DC@���>����lE�u��>g�-�&0�>m΁�~��x'H@K0�>?�g��e��,\?�D��"�>]ڃ��ܾ��C@�q�>����x�6 �>�3"����>�Rt���	��D@]��>m�=��E��>�:�r��>�qw�7Pྲ�C@��>b���d]~�6�?��>�X-�>PZu������C@[��>��2�jP�����>��;�$2�>)�����@@q��>$Џ�I4+�r��>�G�@�>#����:��E@�>Q����1�z4�>��E�ơ�>�+����ѾDXB@�b�>�Q-<mA-��O?�n+�@�>{4�������YC@�/�>�#�<�ur�X��>����>�ey�X����H@C��>��=��7��	�>À'�c�>�!u��߾��B@��>f]�=�6��� ?7=�<��>�Ⴟe�侦�@@���>��� ����>;�(���>3ӆ�k��G@}��>�'�<-'E���?��o>���;ž�(?����~bM=������>�.�?��O>I��+���o�?���m>D���<�>��?Er>)�����Mq?\Ϟ�k�=�����>�q�?蘭>�Z�	�����&?�Z����2>�w�`~�>C̝?��>%�1�����=�
?�����=��4Ԗ>��?�֕>4��~���?*i���
5>���(�>A��?��>A�;������?x���o=����W�>��?��>�͙�eO���!?�#�� V>Z���Ӭ>�0�?Wk>�j��龿�$?�̔��>��� u�>7f�?���>^�ͽ�sƾ�?~ߟ��#J>��Ō�>q�?��>E�G�/(����?N��pӣ=R9��C�>=��?_�Q>+�>����Ϣ3?,̞����=������>�Ǔ?p5�>��ܽ~Ͼ��?\Ó�ZI�=Ʋ	��>uG�?�݊>q�B�mHþ��?�����GF>ؕ	�M�>�'�?V��>Am�u�����"?�k��#�=����>�ē?���>{,��E��۷%?^؝��:">��oO�>7;�?��p>����K(�?<?Y�����?�e6�~�¾��)>��d>$���1|?��!?4�
���?�v5�S�A��>�Pn>Dʯ����?l�?��a?�.5�~��شz>�D>�~����?��8?���m�	?Ep<��g̾� �>i�>д��	@�?�D&?��A  ?��<����WQ>��@>צ����?z{?��a�?3�=��=���>R�>����G�y?��?8l���?Y�=����:>لk>Ѵ��{�?n?��⾟3?�$4�n���W�>�̔>����-�z?<m(?�L��b?-69��z� �\>)א>4s����?(�#?���Ƥ?��=� }�M�.>��>� ����?`6?����?w.;�����ġ>�T>ޠ��oJ�?B'?�-�l?�>�{Ѿݶ�>���>�֭�_A�?r�?����!��>�<������`>�l�>�����{?
�+?�N澎?'�9��ؾ�c�>,]>l�����}?��)?߶�+Z�>C�8�
�ɾ'��>�hJ>*X����{?�?�#���?��5��������>6�O��$�> Ag=�n?�{&?���Ɉ�>�m ?_�����O�.C�>ܤ�=f9N?��?g��:+�>��? @���J��s�>���pn?�.?ٙ�����>�+?n���T�`��	�>j�X_Z?A4?_v���;?^b*?����N�|��>�4���]?m�?{����>�6?���&NH���?�Kϼ�zN?,?�}��lR?�b&?��Z�W��m�>�Ѡ<%t?I�?�=��(��>|�B?V����G��a�>$�=��x?�Z%?���i�>(?h��@�R�\r�>T=x�e?_�?x�����>�l9?�f
�]�dI�>�}��fT?s�0?kj�K!�>�77?���e��
�>.��=�A_?i#*?k�����>�Q;?�7��AX����>�e�=$Au?��+?m<��n ?d�6?�����^�X?�J<�xU?w�#?������?:%*?\���Z�p�~A�>H��\�Q?�� ?��(�>��,?�o�Kq�Z�>ق��9m?�(?����� ?e;?�a��p��;�>�<�;��O?;(,?������>V'?�jﾢ�>A�>}���g��?�JX>���������m�??.0�>�;�>_'���?~֍>�)��)�����+�7�?�;q>�ϛ>�ԍ�=Z�?�L�>q����;�e��6<?�|�>[`�>ÂE��h�?�eo>�X�����������-?�n�>��t>�˞�Ք�?HD^>�����	�2��]z7?]>�.�>:���Wg�?<nk>V��%������o=?�X�>��>��o�a/�?j�>�����!���,�;]?�\�>ˎ>�F?�'�?4yS>�c��t��u'
��7?tB�>��}>Q�R�c�?6�>M��2U#�'f`�k�2?s^>�ȴ>;���oa�?0_�>+���
u�����,'?ޥ�>�r�>��H��+�?b��>�2��. �����?�)?��S>%L�>;Q3�/��?���>����a����??�|> 7�>o�N����?��>u<���>� r��*?떼>��l>������?zg�>7b�� ��tr���@?�L�>}�>�	b�#��?(�>�ƃ�^e ��b���,?�]�>,�>�B^�5�?�z�>M3����J�K-?t����>�8����}GV�j�ǿy�"����u�!��<����>=U���ֻs\M��<����,����ߵ"��:4�D�?��T��Ԗ=��,�F,ǿ�'�,;���������?UI:�ߦP���޽�Ͽ-�'��W¾ɜ!�T���7�>m@`��Ꮍ�:�P�Ŀ��8�L�Ǿ��!��m�W\?�H��[�;���ϿN��O�����f��Ӧ�>�7��-�<*&��YĿy��T�ξo��l(���?�:Z�p^�<��#���ƿ�&�D���+\!�
 =�
)�>�&[��VL�M�����Ͽ�,�`�ž7]$��������>��M�j쭽1z����˿��)�����u�"�����L�?,\�|d�<��)�����]>�����!��L���&?��A�� m����~�ȿ�:�P�Ӿc��y�ٽ�=?cqW����;μ�п�Q � xܾ] �J����?�8_��m��ge��ؿ�K�9��j����$�H�D?	<�.F�������ǿ��!�ދ����#����oQ�>U�B���=���8�пW��Ī־���J7忋p6?�����J�>ʥ��8�S>#��>���=�R�=�Gۿѹ"?Ɍ�q��>|z���c>�ņ>4Z>λT> b�,J?%��%O�>,0���xy>9D�>߽�=5z)>>�ܿC�8?宽��>���șR>3��>n�&=?�>����:?�DT���>�*��XXk>3(�>Z>Q
!>ؚ�=6?�Z���?�>f���(1�>�m�>1�>�_>l9��'?-RU�gN�>RC��hDs>scV>+�=�+�=L3���?z���+�>U����%{>7wT> A>-�=�1�!=1?��E��>�K���}>��I>���=��9>B��+�?��$��ћ>� ��@�m>��T>�W,=1�'>���e�?�������>�X���?>�U�>�+>Yq>�ۿT� ?ݨ[���>T����->�Q�>��
=)go>���ߴ)?q&ս?U�>����dS>齄>��a=}�>0ܿ��7?��-|�>����22~>�r�>YY�=M��=�jݿ`*?���Ԭ>�؞�N:)>��>�S�=��'>t�ݿ�	'?�Δ���>׵��\ɑ>#��>�v�=��=%ç<���>2�?���;��B�>�xþs�i@ݽ�G㾽���>�_�>�� �Ѿ�S�>#����f@�:�d�F�>s	�>�Z�L�¾�й>�����7j@���?>
=d9�>�D�>x���"^���z�>]̏���e@|��Mz��.��>��?;^��Bʾ*�>�����j@�G�}��\�>*?|yݽ�����>WԮ�!�j@E׾u4ʽ�X�>.=?{���̵��T�>�뇾��d@�ھ��F<0�?��>0���y飾���>�k��-Oc@Aw����<?��>C|�>C�P�V�ʾ^��>cJ���k@����Y��2J�>��?ˣ������>��Ǿ��h@����!�/=��>��?�V^�2�Ӿ���>AI���xj@O��q��d��>k��>*���|ƾ�&�>���~k@���]�m�$8�>���>%�	��������>{
����k@
�����L�>I-?�(*����:q�>E`����a@��龪��;&V�>5��>=!��Sپ�ڧ>����h@{d۾�16=0	�>O��>Q|<x�����>�E��9�e@ {�sv�?��ڽ
Ws>�HI��L'�m?�jb>��$=�:�?�W�.��>R4鿦Փ��m0��j?
]>�<>��?U�C��
s>����O���3�4�?NgE>��.>�Ʊ?s�`�e>jJ�,=��������>.�>�0>�ճ?	��;#>�O�\I���E����>�Xo>6
=�2�?�r���L>
��H=���_5����>�yu>�e�=�i�?�h���e�>ܖ��0���H�.�T{?~�0>b��=���?}�*�<�> L��G�����>�?�@�>�}�=#\�?����;>&��揿f����?��>�H�=#�?��T�P>>z忞���&��Q+�>�n�>Q��=��?w'��NN>���<���4���?|'8><k>�H�?#�#��[>�������(��)?�BK>�h=G�?�k5��`f>����6���
�%�f-?$�0>��=��?�Y���9�>��5��*�%�ځ?��S>��>� �?�
�����>8F�����n�dZ ?�Nw>��/>��?��*���>2R��R��X�/�|�?r)1>��s=�y�>Uk�?��І�>�)���:�z�b�.?_o��c�>kL�?4P�Ԥ>��־S5þ����:�?�i���>e��?Y�Խ�C>�����n��:h?+BĿ$�>���?1�"�0>�Jþ�>˾�c��`>6?f����>	�?�7����>/Sþ��޾}��J�'?c�¿���>��?�G(��#r>a��[]���C��K#?�诿�ϣ>?��?����إ>y ʾ��Ӿof���/?�*¿�	�>yx�?����V=>�|վ%)ɾ0Ӆ��?�r����~>�Է?��Y��q>idپ}����Ŋ�Dd:?�����>�?�;μr�x>���������/1?-���k��>���?��'�ۛ>d5�������ڜ#?�`����>ѻ?�(��;M>��ھ�󷾺�{�b�?9���q��>�<�?�>��*��>�LǾ��Ӿ,����*?	vÿ��>;�?�#�*�b>3gľ��������"r#?55ÿ_ӟ>Y��?��0��L�>+�ھE� ����7?	;ÿy��>�l�?]9�P�[>�߾o�;�r���98?o��UT�>���K���%����>��������>�O��?����.��坽��>�O�:�	�ȶ�>�[q�o#�>Xh����._�uʳ>Ǟ���]�>2}����>�M�ˠ�#��<׎�>�!�h�� �>ɥ���?�5����j$;;H�>�7�t��>"��\a?�m��|��Cz��>��������>��6���>g�gն�������>#��kn�b
�>u�7�>[��_Oܾ�;���>/�������>@C^�� �>1��������B=��>�9��"����>)��i
?�k޾� Ծ����V�>������W�>�&��pS?L�H��(ׁ��P�>�h�h^�n�>c+�q��>��S�Ͼ�75�͌�>����5��>�@��l�>�
��rʾ0�5�>u��os���>^Z�%�>��C=���1��i�>g��z���>��L�=��>0X�W�쾫y}=K��>�������>JJ��h�>���b�E��<g@�>�q�����T�>#k���J�W])?����_Ͼ�N�>��>�k���!>��=q�D�y?~z��������>(��>>ė��Q>z�=��H�]b!?T�e�L����{�>���>p�����R>T�=�I��T?��罔%Ⱦ���>�.�>����I�=z��=uH�-?���*P�����>�>�*%����=b=��M�o�'?h��D������>�L�>Z%��x�'>�G>g�M��O ?V�T�����gp�>��>w�4��T>n�]>E�I��
?NZὕ����>��>#O+����=�Y>3�J�c�?t���᯾���>���>�k|�4%>�>!�L�� ?�Oֽ>C��=��>�>�>q;|�Y�=F4	>�cI���?���q�����>��>#��L9>.H�=�M��t?TzO��Τ�y)�>i�>%w��
�=��M>��L���?]�l�R����t�>���>2W����U> r^>/�N��d0?���".�����>���>��z�չ�=�!l={�F���?bV0�V]ɾ�>���>�+;�\�(>_��=�nJ�9?�`�����+\�>���>�꘾%��=���=��I@�����$>Yq ?oQоV�`��<3�[?��>;�C@�>�
�>�+*?%�ھ�����/�ytL?�D ?�jD@���E�>o�?�a���& ��"�=׿L?0�	?��E@��ᾊv�>��?���������=��H?�a	?��@@=|Ҿ�rZ>��?1Dܾ�)����=Ͽ^?�>��H@ ��1�>�0?sҾ����bp<�}b?ơ?W�F@�����_�>U�?O���_��4�=WY?�;�>J@K�̾?�M>yS?���sm�y_U=��P?�o?�H@#¾࿃>�?�H��ٹ���<�a?j��>��D@�X׾0r�>�k$?-�3����;A�=?
�?}I@�Eվ
Zb>]�-?X��������=l??U7�>��H@Ijʾ��,>�?���Q�W6/��4`?V�>��E@oO�.-R>3$?G�Ǿ���9�1=q�C?���>5�D@�o����J>��4?N����~�=*K?:]�>��G@�Ͼ��3>/�,?k_����=s d?Ɣ�>g�E@y�侰^�>e(?3!�Sm��,�=g(`?���>a�>�P��'��٪�?�,z?�]���A�?Е�>�ޔ=�x�>�����F�XH@��m?��9m�?�ͮ>/�=���>{թ�򴜾���?�~?�m�s��?-�{>��=q��>�pf��`W�S��?0[~?�|���?��r>�-�=5�>#���)s�c��?�-z?����9�?&��>b��=��>5����/�� @gy?Op��5�?�É>B�S>b�>4k�B㢾��?��?Cs�����?��>���=���>��󚈾���?�r?*#^�"�?��>^1�=/�>��t�H������?��y?�ⷾ�:�?̞�>Y��={:�>UxK��yQ��m�?�݂?>Z���?x�>xL>���>5�@�J����?�vo?�\��O#�?�?�>�E>��>+zT����\@'Lz?�[���J�?���><�.>�>�>�����@\�1��?-Ny?vm���?$��>ɒ�=��>�$轓�?��D�?u��?�
�����?Ⅼ><�A>�>����H+����?��n?+���u��?F�>53�=w��>S`�
앾�@@M�?�T�+`�?���>�W>PK4'f �   �  PK                      archive/data/1FB  �C^�婷<�E��bF��#��v?���ż�:<oao��4�T!Ҽ�uڼc��<��k�I�$ѩ=��<�=�PO<��k=�q���<Zc�;a��=�nu=�,=f)	=�� =�y��.u=��`=tVG�ߡ��(�f=mN��l;�4�<��W=NVH=�=�5���C�dL��%^���:o�=��:���O�f���7�u�=��=95W=Q�/��=�a���	<�=Z������M��bG�<=RK�vRt=�ď�PK��Yd      PK                     C archive/data/10FB? ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZʏ@_
w@Sm�@���@PK����      PK                     4 archive/data/2FB0 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZF��oYe=�Tf>h��lܗ��{�>�O�����>K�>
,	�ՄG>���>�M�=��>cTX���ѽT��X��>�����a���������?JX�=n��<��>�5J��ER=k %�с?f�a>|��>Xv�>`$>��b>�[�>~�U�<෎>o}>�{>�%n>6?��=��?�2"=t��>�;>lp����>�d&=r�=���>;��>�2>G��>l"�<0�����Q�>t�=`��=`\>r�2>L�>PK
��2      PK                      archive/data/3FB  ��=�@��g�<XQ9�g=^c!>�e�D+B>3�=� ,�vZ���[���CA��Y�;�a�tÌ<j�<r�:��Sh=�-O��&���:�@�=cv=v=E>��=�;>=)R<7�v�
���R>y4#>�����~J1��u��3V=��=�{�o���aث��6����N�g�.����x.>e�=2�����\���<��<$e��Z���n=^�!�����<�Z�<u��uK���f��3t>PKY��      PK                      archive/data/4FB  ��Cڷ�økD�	^�+?��D(O�D�HD�n!D���C�l�E2�B��(C��&��#5D�f�D�A'D������D0�B�#�C��D�@�D*�#D\!CŻ�D~B�C,�I�t����^���u�E��Dgu1D�<�B�Ge�j�ē	BD�0�B艎D>0TÓ(*���ĨP��2�I�e������/4DTwj���
å���}/D�!�����Ù�K�jUuC[������uD�����®�9��<���.Dt�zDPK��c4      PK                      archive/data/5FB  J�2J@��I/jJ$A�J�`J�Z�IdDvJ�M�I��pJ��%J��I׃rI8JTk�I&J�uhJ��sJpI"��I���IhƌI�	�I��I��-J}��I��RJ
��I"{I�˭Iv�J5J���I�JVI�6JR�tJ�}�J��PJ��I�&VJ&��I��Ij�FJ~��I���I1�VI��DJw1�I�GbJ��J�	�I�#JC3 J�9
J���IL�I$J�\IF6_J5�xI���I���I���I��I$�IPK[o;      PK                      archive/data/6FB       PKƵ��      PK                     < archive/data/7FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ���D̾:�9�`�?�վ;d���#��L�*<6fQ�d�����E�H?�cF��cľ�3��4�[w'?/=>	�c>J�?[�A>�<ý�V�)?7��<+�.>as�>+S�> Ω�:ʠ������=�"� ɪ;����=�=��v����<�>��v&>�ɾ�b��3z�_]��1鹾zZ�>�ƺ��TD����n�I�D>�������J��
�>v=6����\G? Z>����zx=��= �
�WE��>�����]��$$M=R ���?={e�>
�?S>�������<_d�>���>���>�d&<&c�?�@y���A�C����=�;%9�h6g�MCj�Oؾx�3�܃��y������YP��+��奾���� �=� ̼\�v=�j���J�W����I�rQӽ��̟�<��>�?��&?�;?L� ?��,�$�ɾ1^�;&5�>�艿���Mg�=�b?BbȾ{�i��?+��j��(�`��P��6վy��=���V��>sL>Zs2>,m�>�엿]>,ql?�'��?J����?}��Kz>����z?�3�L�?�����xg>g��?�b���*=7�q>W�⾩٠��KU��r�>׽�W�>�N�z�)�E�Y?h.h>NR=���A��վ0]]�t���T4����Q�asS?��m�.ڕ>?���[�8\�>19� ���H�q>����l�$�a����S���>8�n��ؾ{�5?L��=�jc��(w>/�>�W�=��p=��?�1�>�^�+�@>��2�[�=HP=�%k>\�*�Z�{>��>e%?s�.>��?��8���a=���>��x�&%���H���,=/�>e�4>puN>�Z�$�=���
ܠ>'���%@�A�Ͻ��N>g�;�0yr>�.J>I@*>�l>4�?I�2��0�=�\���4�����xϼ+��p%>�ξ{�N;�"���(�����>��>�6м"D�X�ѽ�B?�р�)�'���ր�>\\����i=��� ?U��;�� #%<?�kYr�6�6��B���&���ӽ	���M�c��=��,��� �>�{���׾{�>Ks8�*xL?w��=� ?�L�> ��?�ǻa��>@��W�?���p7�>K��jr�>K���z��s�̵����/�r�6>�j>� �>����2?�n�>���<��,��>�Ϫ>r��?<�>$�>#�>t�k>u��>��>��>hE�F>U����>$F@=��ľ�k�YR"�N�!������W�=�T?�'�>a�>��>�~%?�D?��>R3��q;=R�?H"r?��q>;b����<�x�=���>�'�m�$���>�E�>�.��آ�OC>	/_>g�G�URb�J��>�V�>�C����>��*?��>�=f�>I�?��&��U/�@tm���=�����޾U�&��Tξ�F������x�����V�}��b?��9�b˽�5������M���W��<2S޾
w��)�"��>~��>�4>(X���H>�㚿�[K��+]=[Vݾ�����>�Mϻi�@���:���=��ܾ����=�[>p׏>���=B�G�-▾�o���}��޾�9T�/FL�.)��Ô��v�=�в���:����>U�i>��>Є>�7���;��S߾��7=A���f#q��"^��R���N>k��f�5��rm��==��>��>Jc�>�q�>�&;�A�>G�>�$�=&�=�(�>#5#�=O
?�C]>��ܽy��>J?S�"���i��k����7�Gܓ�X����ھ�2>qپ-޾W�;�,�
>x}��a���.t�'��>�!q?<ɫ��L���>���=��>XR?�T�>�*D>��>���>�=�,>��>>��>8��g)��������?o,d<Uj%��9j?2B�>/?�*>6U?= =U4μ_I�?��>��;�y�>�[����R�w�`�-���3�O��&��8���4������{��Iʾ	T���ľ�/���=�9ӽx�H>����Jtz>��������.`���V�T{��ʘ��V~��p�>��پ~��=�%/����=n�ӽ5 ?bˎ=�~�#�>t�#a�>��,�``��"���gU>��
�+��������C���_��1��>�3s�
�e>�K$��]��t>'a�>��d>�)�=��=Cφ>b�
>v�� �?��<?�E�
A����i��F���?(�C?٬����%�S?I�R>Z���X��>�
?�3?�Z�v�?��1=����?��>I�?�G�<ó��#�o@-�li�M7f>����6��v���I|r��`�=����j>�,?:��=�݁>���]ݾ[ٛ��7���qu=M����ۣ�OL��Iν���������Ⱦڽ*>�@@?�j�=�*U��>�t��6}�<m�>[�b�{�3������>4�=+YD�N@Z�2�g>fMH>>>��T��>iۆ>��?�)?�M��;a?Ī?����&��:�>��=5��>A��c�=�������8l?��p=�<>�&?>�	?K�?8J'?M�?jLR�@`�=A��>�`�?��<9s��*�����pH�<iu�>�V;?�%ξ�ن>_}���\~>;]h�}޽^$?%5�?��g>0�Y��>�m�>����SÏ>�Z�>�l�>�R,�oGM?qG?x�?�M�>�?H�3?��c?�H?y��?4��?��?�	x?;�-��'$?��[=?*q?$&쾈>�>7��>5ڧ?�`Ⱦ?���='s�?��>|�>=ɨ�^?�{��)��)�>.	U����n޷>C'?ʄ4=_�=@<�=e�=���=[�<�!u�G�=V"�������0�>`�ƽ��W���&?� �=���9��=y4�>��>����>�0d����> �<[E�== ��{�qQɾ�4<����s�ʾPd����^>y�y<�(���fb����M/>��>��!���3?�ʵ��:���w�R�M�c@���>/���y�A�f3�>Y[�> ??�� ��z��\>�� ����=jt=I���H��n���P�GI>:&ɽ$���B����>%/=�K�IU�=�?X�8��C�Z8�\A����F��Z?=�H�w�m?�G=ς�?Ի��ܾ_?��T���?����(?�S�>B�?%�*���W�-?��? O���H>7:�>ݿ����	�c8�����=�҂�wn>�=!>�s2=Cj���2D?��=Ӗi�{��bO�>�(F?Q�1?�[��yd>k�r>7�8?�/��J7>q�ý�O��[]��p?�,>�����f�{�&>���>�����S<����>Ⱦ=��>S;?2�=�����6n�NW�>F$�>�㗿�g���.?F:�=7>o���>`��l
}?G>�Ձ�*�-���b>��k?-?*dv�$�=�x�]�>�T�>����y>�3?<�>r~r������>�"��3?U�??��>�'A?䴀?f���?���??MD%����?B{W?�>�h�>>�>���|��z̟�N�c>���c��׮?�0 >�hپ��u>@?�>�_�B<I>�=8=�e>�q� /���a�KL佋B>�˩��Ð�A_�1w?DK��ZZ�>�k��I�=��?D8�>���>���>Q���|�=[�%<k`��Wa���51>���������>;U�����K1��վ���6O��\w
>M��t�?%d�=&�?��C�z>���>�xO=0����2M>�@�>�>
�߾-(O�CR���y)�S����*��T��4#�>���[,>���</�Q>��=#�>�]¾��>�W>~��X�m��bF�݄B>(';�G�5�����p�i���C��=}��$?1T5��	�>2g��&>�;��P�>��;ji&?�&?ӂ?�N�>	��=+Nx? W2��Ͳ<jBp�.�m;R���Wxȼ��� >Ndھ�� f��!��MV�D���̠�4%<�z���!���ֵ��'n��7��Bƺy׍��e�>�^5��O�>Lv��8��>���_�=�;:?��?]7�>��Z�!Q$��v���/Ⱦ��p���?�ʣ�yz"����YF>{�?�?Ɂ?�][?˞?;UB��K�>t��>Z��?[�C?/so>��^��	K<�}����l[�RQ���?_݆��`?�.��(H��(n�F��"�6>޾`�2�k�1?��>`��;�ؐ?H�>�����>�q����!C�>-� >ڼ�>g�w��1?R�?l�{��8��m�>?�?����H���p�`s�� *�3���e���0�ϵ?S�Ͼ�tV�if�=O(��S>n&Ҿ.)	?�l�?�?d������$��D>��Ǿ�Aؾ3��*T��I��V2ھ5n�����>e*>��M���5�������ބ�=$���A1	��J����J�H�����iM������*��E�>K�(?��%?_bB?<�V?�:�>�־6W?`�r�㠵����}����> 陾"�2�M�s>��=Q]��ج��I#�s��/��>��B��M�D>C��=�=<���鴾����Æ�5�
�;@�>ݫ3=��F����i�$�j�?�>?ߕ�?�W�?�?�>����6l�<�R= O��2ߌ���þ��?f���WX�Q��|��>{X���q������H����y?|���W�?>^>\qB�S+F>j��>?�?��\?�	�K
&?���>Ґ=���Iԕ�!<�"4ԾEѽ�UK>ZSN�3���U_��"�>��?զl?tG�>3`����<�<F�Deӽ�y?���?�O�>��p>m<�>���?�?۾HZa�.9I��=����@��7�>h~�>�g�����'ӗ�MOz=Fu�;K%�>�W>�f1>,#r���
�W?̓D?O�?OX�:,z?oK4?վ�>�M��?����<8�7�?L�g?�y�;���=���=Ys?	[����9�+��&J�`��)��>�p?q�"�KAv>-H�=H.�?B����4|�|�����?겾Z}+>��-?%2�?����sJ�OT*?��n='�?(B޾a`���Ď?
�=�ڠ>�v,?K�ӿ����wA��Ƙ�^��ǿ?�T����q�.�5��܈=�+>]?�ؾ��"?��P?�o+>X�O��F$�S��>��������,5�) �����֝�2(����>�G�>�ܸ���۾��쾔Zs>U���t-�>Y�?#�?��=뺐�\�9>L�����[?#��>�>��%K���t?&nL?�۾b�`���޽�-��＿>��$(�>�%l>fF?a����վD?�^�>z^T?PB+��ĕ?I��?�!
�8�L��y��P�c?ʧX?�̽��g��*Y��ہ?ӻ����O�[��ȅ�>[�K��7�&m���Ѫ?�9���Z�Qѡ=P7?z��?��q?�9N?3�_?�mc�9Y�a�����>��ʽ���>?j����e>pL꽁�'���46���m?�KO��L�?ys��!��Xb<���˽�-#����m���i�i)�>���Z*��/������f>5������R�ҾmW���A?��Z�V��=����- ��� ھ5�þ�ԩ?�{�?X͍?��h?�8�ۄ���>`>�ht�X�>�Ad�S�4?�g�^ZE�l�=��ľˣ ?o;?mZ�?�[�?R�>6�[=k���x�ؾeW�>=C�<����'.\;�Vѽ-<T�����u�>�% >L������<�'?�>5��Y���-V�#S��,�>�t�<��x�d��ET>��׾�¿���l�ּ������L��&dE�M��=5:F>�#h��z0�`�&�_���O[��������`�%�����(�&/A?��>��>O�>�v?�X�Q�
=�/��R.?/)�>���?��>�?	�%?��Z?�� ��6���ؐ�W1����r��O��-��>�p�0�t?h=)?F���^
?n\��ݪG?���?[e�?�vA����B�X��K��G<@��5�bv�� ���x=������C�E�پn���?>�HD�����L=���>�[:=�L7�k(�>�Փ=���^�>�=k���;ɾ�B�g
I��7Ͻ��W��^�_>��>!�S��=�S��hl��<J��/��>y�>��LM?�M?E�>�F��<;?�_�N>Ap�>�vg<@�Z=�2u?UT>��8?p�U�2ѾO*%��7�?_''?5?�հ>f��?�k
?=i���4>�*���E�W/�Wnݾ>t�=�p~?��
� ��\Yq���/?�ti�z?�qB?�$���?Zg�F3?:�S>�>p�.���B?	P�>���>��L��YA�>'d��|*�>�`�D����>�T+?�}X?i
q?�w?���?����W��|:��s�D��<7N<�s�<�>4�N$�S�����٧���?��>�-�>���"��=M�]���>���?Z�ҾDw>*Q�=a��?�T��1��q'�f7�?�g���'�=�?BG+?�R�we>�?G�[>��t����?��4?:Y�?>`s���]?N��?p?^���l3���ھ��>�F?aa=�:��֑��- �?��?�̿?�xA?�?��[?�Ē?�>��>���ﾆ�Q��A��F�#>��X�z?t �+��>V�_?�&�>������a?,Z#?�<����'�M��Ә��/�3_U>g��;
�n�z���Ra?��P?g�N?,� ?c�>z�>.��>�O�>�@0?�T�?�{?�	?b���fTľv��>��>-W����=��>=I ?��p��l>�?��s?x$ҿ+O����ÿ2�z?�"l�G1�=F�9>
�@��2���eL>zj!>��v<I��=���&h9�Z���5�=A7>�������rҾ���z���P�>8^�>���о���>�O?�C�?+.>�-?Fo�>1�<��_A?񩘾�<>< �>9��>Ԭ���^@�#��׾�AF����>!�*��R%<��?6�2?��\?_)?���m���Z7���]��ma=�>�d�<W�>�zU	?�
�<��?��(���)>�^M?Y��Yu����>�����SC�X[��Nv8>�4>r5?=[���
Ƽ�??G����K���#?ᄻ>�� ��P1>+ſϪ���>��Ѿ�O��'FZ���P?u��K������<�+?7kL?��п#�%?���?PG�<�*�>eMt��ͷ=t�v?��?-�u>D�]=�7
�X�\�m43=�N���4U?�؁�O������ℯ>`�[��E�=��,>�����ٵ�RX`=���%��?S֌���W?�E?`�)?-�z�y���KƜ="t�>�1�xU����>3ʥ��h,�F ?���ld�>����-ݠ?��>���>]���N�k�og�!������>T
����z�(SS�q�P>l��>�#�Θ>1��sUľ=�B>H�>?�?���NtQ�(��bc�>���=�`?U�K>�7��M�I��>�,t�B��>�y�?V�g?�8�?U?�x/?��?�L��uř���콕Q�a&�?��?7l?f����j?�H�>�*˾����>�T#>(���4����ؾ{4���C�>O���K��YG?��~>ɢ>� >ū	>"U�=�S����=�T?�]B?�$/>݋���>܆=���>�����-���a����
���Q�/�ž)�ξF�}=���= �?��L?}j?}FY?��|�d����<P�J�F�$6g>�ݻ?V]��͈���}�i�?`�D��� �n�оpq�>�o�Po�>�1�=!�>�Xa���8?�H����?+q����^�����2� ���mcοv�������~<�6-=�,�=a婽��=Lɾd��>��>�>���>��y�+5�dؾd?�Im���Ծ����O�~ɓ�m��.}�=��>#�0�Eb��g����>��
���F��3�?G�?�T�=r�>^�>F������>;ܝ>�h;������>�76?UP���m���qҽ� ?F?��Sy�E:���o>
;��y羯����?Qz�=�-�����?G�G��㧿rg��ei�?"�#?n��X�87;�>�~ɿŻ,��k?kl�>�}?D�ƾ*�w>h��> y��F��{��� =�ؤ>c���X��>Q�L?-�o>4�M>�%i>�ʮ?�lj?W�?��'?�<G)��_�u>6 ?>�*R��d������[�>�?�Ӿ��=?�������-<�����>�N�>H0�>JW=,�=(�>�/?*?�U�>+r���ˇ>+�c?����&'>�w^�����p3�����=0u�>w
~>ؕy={�(���$8���^�]�$������蓾n����4X��%��p�>9�I��=��{?�I?�>mp>@{&���?��>�ӏ>�� ?�'?*��?KRS���:��͛�Ù?��޾^������ɑ&?r�>���>xG���->�J�������#>2� �m	��Rοmi��r�.>���=��>��F���>�:t>X��>��>3ϐ��[�Z�����?Ԁ�������*����>�c�Y`f������q?y5<����B����ڽ�nq>�$q>���>�Ȋ�5��>�v)��e\>w~��J���������c��X>�s������I�$�t[�>p�����=<u>�C�>�R�>.6üm@>:�#?]x(��G����m?�!���k.�񗃿psT>!C�>��$?Q�T��:A�~/:>���>��ɾC����Y�?'\?��=�>b1�>j�H尾,k{>�>����P����M+^���:?�і��;�6*>��>�BY?+��������=�)?�[���m���>�.?g_r���׺$�!>�S¾@Tz��P��ھ��Ծ�ϳ�T揿R�p�[��'��Z@>��=�ξ�iN��R�2>�?���> ܙ=!��>9�??�^>i�F��?�u>��->�H�?0��>��"?(�o?[�y?�qv?�HB��l��)m=a]?po`=�Q>�>�m>n]������6�E�>�EҽS��>�b�g,?��ž4Q?�Ĵ��5T�z�j?���>/eC?�	����>���>(��>�o�>X?p>ŪD?�!��{
��3/�LZB=�?��V>'ݾO3k?�v�>?"���Y�?�3�>Zqj��m����'R?�(��t �4
L=E�?�`�E
վQ&����@��m<��U�'j�@TJ��ٸ�����o����Ӿ�Ɵ����?W����r��L=���>x,k=�1%��/�Q?o�e? ��>H�E��fl>4凿���?ꜣ�aW��񴘽��<O>m�/>��8�8Z��b�?��-����Z�·[�^�?L±<�і�7�	����x��?�[^?mhT���?�=��̗?��#��h��>
;��=X����>�5&���? "7��]>ف���vZ>�
���YV�O�>Om��}(㽟�7�k�>��S��c�>j�B?�܋?ma�?�K#��������?8i��%NH�a�<8pL>���7����M�c�
���ܾw�׾bK��D�-?a��=����#����>�g1>t	3�7�a�)P�>�
�x�?	I >���=P�-?d�?�J?fg���-��o��&������D?�������?�>�<B?ym#>��C>�d?�4�>���>�L�<Ι�����\�������>��?�Kh�_k?e#�q�p?�O�>��u?-D?�">��>�+.>��佺�=��j���x`�=#�?���=C�<}!?�U&?�դ<��>�Z?/��>j8z?�#�>��>���<PxH?�3?D>l�=2=����$���� @I�U���H�={�]����|o�j�w�E�F��n?
t��Qq��gt���߽�ُ>�"�=�r��PY��H?�_��lS��,�>�fA>��=�"?I{�>9��?�d�?��>-瞾w�H�.��>~�>7Ͼ�E��{վ��S���?���R%"����E(>+��>��>����B���I/��v��b.�>	�+�>��Us�ʿ�L!?�L>�?>(�?��/����)d'����>S�����h� �d�����>��>�#�>�QM>�0L?�3?�|�Ӷ?+N?Ȥ>Eq���L�L׋>vM��üV�L>�V3?��=�<�>�2?L��!��>㰘��'�>������c�>Z?2��>�D�<-�`>%�>��.=#>dn��5�>�頾x{�ʖ齉.�>%��zf+?X4?w��<卷��9�>_�s=�m1?r�-�I�r�&6���Ӿ���y>�#����z�y��?L��>��^?��-?v��?\��?a�t?��t���)>uj�>Yx���?�n���=(>�O�������Mj��eG�	@v����>qh ?�=���6�m>��?S�y?I�?s|��G��f�����d?�~��U�ξ��;�%��=��̽7����U���L?�ZC?.l;Y��3.^��5>�В>��?_��>S^����}�Y>#!��jt�أ0=H..?�2?�㔾_k�>��'?R#�O�Ǽ��>��>�΂��t��x?kε?}㔿�&����>і��H薿�Ծ�X5��Zx�@4�����?*:�������?��>9z�?��e��c�P{/�s���A���Y���n�;���F��DP�=�C>�=]�)�O?�?AZ ?�־je����]>�L?�$��������5~˾U��*�+����=���>�߽z4/?�MZ>�>D�t>d�?�{�>=e,?�O�=1��?��?(��?��	�N��O�!�u?��4�����?�>Gi�?D@\?����X?>n?�o8?y䟿�`�?F�a9��TX��Z��>F�ؾ��|�ѽ�d?�Y >��)�6��>��?[n�>6�j>�s¾ZH>��=>����꒾'	�?�D��G�>�\�N'N>�?}3H?�HA�-��>-�?��!�* �>�0��0�<?i�
��
>���1?����n�>���S��b��?�
R�������>q�$?��7?��9?�>l�#�Ĉ>i�%?��O�
?���>�QK�����E�=��q���_��q��
.�=����Q��Z�U3��NR�����B����=I^o?�;b�m
=�>	?�-J������1�f���N��>J��>�\�����Љ�袭?�♾������>,?(f
>E���<�Ě?�>��w�-G@>$�Z�R	?��?�D��C�K����>�%?>F�l?���!�����k��OϾ�L��D���������پГ�>s#m��f5����>?�h���X��1*>rP�?��,?�о#��;���=��U�R@o�H�]�{߅�#���K����9>���=��B��L��X:��Y$�?`�?D����<>���y	|?P�O��0���W��ܾ���=��+?$	�>a�����E>�d5�GO�>qP���[�)���Ke?��'�U֊��0���cɾ��>��-���X��ؑ���@��ǿ�f����V��)��uK���V?�߾
�I?�+��Ff?�%�?b��>�Ե�EŊ?N�X��	@="�?�.?��۾Q[*�S�>�8?���D��.m�j�MC���.�=K~>r�?ރ�=��y=�*U=eJ>�5>H�y=Z�?�Ј��} ?>�Fg�=�a? �A��1>�<{=y'h�c�`���a>^L������NR>��=���=�<�E���U.=8@?�T?dm =�1�>�=��dI�=�X?`�v?�ss>"�l��l>��=�w �(G����ꦽ�՘>%ү�M�Y���>>�=��q=�|��fv�?˙[?��A?ٕ}�s&�~��.[�=J�=^w(��׏����.u��8�ƾ�?�;��ս˭��y��>��-?�R���~b���P>��={kսz�>%o����>M,ݾ5Jr�y)r��v�=�>�>v0��d�5�?ӧ ?V�㾉*���B?Ce�>ٚ��)�>���>��?�H�?��_?�G?�4#?p�?�>?�<	���	���>3?������?�V�?�=�H�>ֿ��q�?�Џ�;�E�� J��x�&���b`K��ZN?#O����-��'>�cEe?u�I>������>�*Q?G2�����E>�;�Z�Q���� � �J�<�d^\= 
'��Z�W�����Ž�bž}�=�:>�
?=�B?F �;"K�>6�������S?���>��6?�S�=�t2��V������O�
�#���络l]�7@�>�.�>��o���>��>��a�!=؃���F?½&?�]�>�?���>��|?�7>�cI?��Z>�N��LH�LXz��%��"�?�ܽu�>������=݃�>��ڽ1X��u����)ξ$���������c�?�ϻ��&���>FY?��I������>wķ��'��o>ʗ�=��>�R:?>�<��[�3��ʹ�=([z�	v�=:�����<BQ>V	������>l������T����#�=��>��m��>��?>�̉����)�>%h?�?��8?<q ?zF��h�I��K�{�Q�-Y��3��"Ӿa��$a��d7�u#���=��1���RѾ@���,L?��C>��ɾ�|=>�U ?Ǿž�j�d� ?!��o�@�,m<��O�>������>P5=��V>'�F?���d�'>��>��žY�/��6a��2 �BQ�w'�>:\�>5��>{�>N᩿ku�]</�YB?)�{�)m�q�¾����M`?�]=1��=v@پ�=ۙ��>>�4=º�>i)�>k@��徑C�i.��"�˵s��k�>��ľc0�W"�=���>�p>!Ҫ>�^>���&�>�����?�w��c?��5��=�>6����ž���>�>�>�,�����Kx��jG�jύ��y�=R������FɆ�FA��u���>��߾L^�>r��>�Qr=�,�=Ϩ����>I-l��W��8}a?�<�>��8?��5?�i"?�L�>�Ϲ�T�>�??�j���L6��7B���X?�2N��$?nr>7Ͼ�CG>/���
�>y�m�����{�e�=ޫ�>�ۼf�=/xY?A�6�^=P1���$-?��;?�` �^��F��>�Uc��vg>V�>�E?;��+Hi��Խq�?F��>����U0>+>�����S?��m?i�?�cҾ�{?�8"��==\�(m&?5��> }ǽ���;�E���G>ʻ��	M������/���l8�y؏�X�B>�}.?DN�:�ܽ�֕>*Ņ>d�>����v��>�3���н���>���<�I7?o��=�	��(���4ؾT,��fgP??�����>,[�]�3�SN򾌽v�~K<Ű��j�?��t?ﱽ>q��a�>oې��p�=���߈>r���Ǩ>���l����A������j���=�|�<�_O?��K>G�/�'�[���?���=����/ʾ�(g>3�>���=+ɼ�V>��F��0���:=��#��Su>���v2��*���y|�>HN3=��>j��6/w>�����YJ�����bR=��BL�h6���n?�`>��~�\I=� *>X�=������m�>x��=DJ�>{w�<Ĭ>��ӻ�$#R��y�����
>�ν�̹>9���o��=M�"��g�Ӣ,?���>>��?P	Ҿ-%�>`}>A$=A�>��m2�;��>n~���̯��UQ�61?R�?��A?�'X?7�?1w4�]L뾗����>�p�=�n
>�+�>j[S>Ə3�	␿*�O�=p�>���>�H�>�{�>I�@>/
?�~B��M>b�?�Pܾ�F ?�������:�b����2>/+<I;?��>x������(��0�Bn�y0 �}F�=���P|���V��[Q�>�,�>��޽�+þ����
=ָʾ��)�;F�>�7?�ަ>��?��;��r����������!>-�?��?z��oZ�x�u�˯�x��ਗ਼�ײH�(�g>�+?胾:'M>LM�=���6�a?�/�j��>�L/?�����=����6���u�=kF�ǚ"=�!�>C(X���
�|�< ��2y��݊���P��-2���>��I�/��=ˣ�>�*=Mq��ԡ�P'>~o�,�뾛�/>��">�����&������N��0=��6�k��>�>/l!��R�PrT�U��>��>��a�	Z�>�:�>�e�Y��ƛ���s1?B�?h@�>ɋ�>i0�>r�<>�3�?�)?,� ?�=�5���W>�<��C����<>4v�>�bQ���S�u�#�I�B�&�-��/��|?����¾\�y>��#?�7�>���>�fu?�B��ڲP=-���Ҥ#�-2�?���>��5��?�(9��5׾L�b�<�>�$?��\�>8ͼ�o	�I���$1?ĸ:?��v>x!S?C>YƲ=r?]����_Q����>�	?#�>�;�>�I��Fo��˽�Lk�>���>��������K�>?��>�_?kv�:��xh���4?��>��=E'�=�y%?G����b��'>�bE?J�S��,	?s�?�*>"�H���?
z���lP�2�d�9�>�g�?��G�G&G����ݝG�3�<6�>�]?�\?p�e?'��=�1�?���.��F�0=�j?pDO?�;���������@�&��]��D~$?k`��k�?c���Қ=���L�ϩ���VD�I��>�wF>�r?5���%��00:���W�ͩ?3�A?�?L�>�PV?�Z+?<�?���>Em?.�!?��>?�?�J�>Y��>v>��=,�����G?|�?WT�>a���(D?����TϽmyW�#�6>f�>�FN=b��5�a$վ�m���%$���u懾}�A�`Lٽ	\=���%�o��ㇾ��?.j>8;�M"==q�
� �O>��������?����V�[xX��3W?�D�>#��>Y�?In��h��BνB���K�?Z�-��_y>~�{�;�M�,��B��f�=�b_>S'>Q)�>_��>K3���Ӿ}m>���?M�?/#�>��>3?�?��Ƚ�>?x�6��?Y���ý�B��Q����*?_�w;
�>�?8� �)�{<>U���I�6�;?t.þ�����˾��O?�?�W�>ZL�<����)>S=�"a�%~j=���>�*�=5�%�P�'�T)�XH6?�m�=�J���?�(�<v��>�V���B?|���sӔ��6R��4���}�>��$�\Yg?�Ⱦ�8�=��,?bk!��<����=��Co�t��>R);#>d8�"2����?��m��"�x�_b?���?� 	?�(�҂"?�������X�i�cݾ�x�y>�? "��?�g��=�҈�-�!��L?���?G����R���|?�����뮾g��q�n�`@?�^���⇿�i��w|��	I��>h��>�UM����?Oq?�|��
i����k�`�=3.?�K?��	>>}>��I?�ҵ�K�=;I�>�R5?�������k=�<�e�\�m�I)?��R?%�?A&w=N�� ~>a�=��?���<�x>?���=��/?���=)d�0)���=��N��!�>� = ?Iǽ77-�+�>��5��>8�&�z��;�=m�?&s�HHS����>pY�=a�D=~���i?�=�E=��D���þrh���n.��S��B�;I^�[�����=o6�>p0F�g�>�"�=�s��2��|t�>�nh?Q�3?.�/?13%?^�|?�f;]H�=V�>�O�>*�v>��8�Cf�"D\>��'�L�y�\�<��yj=ھG>-��>���>��qM|<7�V?����O�>��>��=���!�=�hE>[�>!Bp�k��e��>-��<�_4��H��稾�L��2�������>�Jw<�Q�=��=�>lHM>��#�խ�>�.ھ�9>�/׼�$9�F�ҿ�
u<���>�#��^|��1>�?��Ӿ�>�+�������:־�L�>�@>�"Q>=Y-?��>�O%?ȶ?�4�>�Z�>�M��)M�>�Q�>o�l=�wx���s����>y]p���>/�>`�=��(�2W���_[�	4�5 ����>����x�>�ƥ�$�M�&�����>�R��8(�=�K��=�?���қZ?�v��d��CE��^���7[���=>�����l[=�>|�?g">)M`>ZE���>oԄ��Y�>$U?ra)?#�?@�s=B|<�Z�?�i =�q��݆>a%��ݾ���u뾛�?{�:>�X�D�>�0޾���>�g;��5�$&��Խ)��HJ?gO�>�v�=La>6�d>��(=��W���?�"���l=���T��m�/>$2�>�辮������>0�����>>�!�G�\;�=o�����
�c>hEӽ�hK?'y���3>��?>�i>�f?�㫽��i��y4?���;t�?�[�>��?s��>�G= �ܽ�Pξ���eC>��>x�>��>Gн	Á��n�1�y���<��P��پ�`=���-�	���>�a?�b]?vS:��]L>򲣾�f�>l��>z�S>�`>s]���Z��}4���w�̙��s��S�c�����V�Ƞ�+����5�b]>�G+��������=W�>���=�p�>��>C��bH�ҵ��Wm����=x��=X^H>�v��$	��Mt���˾�K� �>	,）8�?�K?��C�z+���]:�����v�>��S=��6?��&?�i�>�r�>̍�>�ս��H<��I�G��)��B�n���S��֛<��	�	�>\l�>ȃ8>-�
?ֱ�=f��|}����;�dӾ0���D�����۽L��>g�m��
�>���Β���ѾV@�֮7?{0
?D��=�W�>�>�4�%d�=�j �D�=��ܽ�G��`��X:?;̭�E�q>^" ���>`:��j�L�ka�͂�<G��<��=T���Ɗ> �?U9?��@?_��r?�)f꾧A����>]nl>02�<RL��F�>2>?�?;[�>�?�Q��G��b?�)�>
>�>>ė�kW�>jB��w�k��]�=�|�?g�>G���
�>_���̡/��Z��$������6�8���5>�b>����Ⱦ>�����>Ës>0Q�$�	�N��>�p����f?P�>��>pb���;�Anr������^?�_>�Y��6��u��>�F�Tz�>b���Ʃ1?�6?3��?o-�+�2>s�=N[�>�`=�
��>e�>��?ٜ�������w�)-��F�G�*�Z���2پ����̏�F��>�cG�Av��̷=�?ˉ�=br��tY=#�>�u\���>��>s�+>&p?/�9>*�#���=�2�f�I�� �>^c���3>h�Ⱦ��=�'>���>*/�=���=���>�o1>݀�����Wf���Pp=�z|�7Aj��[t<sqo=������=�k��F�>Tͩ�� ?\�~>�>:����)�a��|��>���=Ɓ�>duI>=��>@������:K����>EǾ>ʗ�ʀ%�R��9���Iъ=�%<�\3���ھb��[N���Q���>��A��Q4�G��>�B�������<NFξ�k����=�q�n�>��=&an<wTc�b��>9A>cSC>�@q�i���\���������=r����#>��>קa���m�s>a�>-Jz>[�->�M�=*�>�K�>{\z��9��7
f�CA�=f�>T��������6��&	��`@?2��>��L?��
?�M>@��=D.�;@�;>�]��̛F<G��>v���0U��<�ݽ�\�<��>�0?W�?8�	?i�˼(�M>��>^c?�=���˽���;�>Ƽ>�����G8��Jo�����_�"��=�i��<$7�A��<��(�5���C=����?�
��H1���&=�%�>�<c?o0ؾ��`�Y>���=y��L����6?e�>�	�?��>G��>��?�L/?��-?�E�>.�����=��=��<>�ߊ��!��	�վ\�=��!?#r�>���>��>i�f>���>��=��M>E�ﾧT0������B�t�]>�/�>w��>���>�p��C�D���8����#�n��zc���k>��`1>l�>ZL�=�+=%`�>\�=$?���>e*���ԑ�W����Ӿ+I?���r��=ȹ�<Y�$?����3
>`;�zw�>���>ӶK�h@�?��W��*�=�Y��
?ܦ�>."�Y̜�-Gy?�K�>��t>IZt>ǧ�>��E>9L�2��<+��>(R0?�_�>�?t^&>��z>�i�>���>T�>'��r�<�p���>��:�>��w�)�U>�]�?�#y>����X>|�t?`?;:�>��P>�$>�d>U7�H>
0{�!�q����6�z�O�l>1/2��� �>1��>�D=��>x<�����@���	�<q��$���S�����^�e��>n��K�>������?�5LO�s��>�ֽ� ?�%?g�;>��>��8�`��>:�۾Ի�>|��>��k=6QҾ��׾ 0����*�/j'�j)�%�a����M���@?�7><~ �=K:�,L辵��*GD?��(?YD?q�<�S��>�%_>�d3�����<w������.���f5��0���)�>�}.?���?T9?@�?��P�pg�>�I�>�X	?�(�৯�{����g��HJ3>?Ks?�n��6p>q+�򺽾ge��)�>��>Վ$?�[=�>�қ�z�w���=����>~7?�u�>,��?ev?)9?i��?~�?�>��_>A�?տ?��a?Xc?R�W?ک(?9SϽ�������l�N?W9��X�=� ?�7�>T6z�x�W��;��/>2�r�H�-��>�Jz>��ȽǙ���G]�#s�=�"�=UW�=�'�=W��>�}»B8����C=�2$= ��>ħ?(c�>%n�=��y�N��>������9�<=*�>=��0��e�?��,+�>��]=M���� ��q�����M�">�ޠ�y�>O�=A��#�w���=r�D�������oF��$��划>�4{>��5��*>a�=�>�$���?R~�����>��L?2�rL:���?�r�k����,�\r���V��q�|����=�PP���-��n�M�ͽ��>9�2?�`�:6n����=�#��Տ�=�>k��ᗾ�@��^�|o��>f~�r	�>�����?7\����	?!Hþ�9�>ڼ>�+H>uw��}?���=��R?1�)��pf>���=<#��M|==4�>&+>>4�>���Vv��덼�w>�i>t
��ɽ1h��ev��-�>�n ���n�SH�=@��?AS?D?"q��|J>p�2>)��>���>ؘ���?�>�,��d�O<����\���pɽ��>.�4?R_Y?�4���y��U:��|��=���&C ��.D�d�޾��a����>�&>lf��ֽf튾Y�\���#�T��>lP�>���ʿ{>Z��=��'�8��>�]>�ս%&>��<!�E�t�>Z���U��?R:��f�1~>�U!>��w>C�u>�G>��.>�^4>NRѾ�Y�<N�w?%=/��>���> e�>�ې����>��?��$?5t�==6?n<�>$.<�����<�����M�1�ݠ���=����<�_C>A�ؾ��־=���[��>N\�>�I߾<衾���?�t��?�������"��;���
�>����H�T=5bL>�e ?Tړ��Z��'��<��>��r>}bd�Y�[<�{�>�_�>�e�>�J��3�I>5�#<�fc���a?$-
>S����O">Ӈ!=��>z���)���H�&J3���L=f��=4�Q����=M�~�FO�u�y�n�?�j�;���>nK���B����U����J��}��X����Y���b�p�,����gU����q����{M�;E�<��y�@�u��������<)��j�h����m���O{�� G>6aվ�)1>�$�hM{=�$���`��H�{��1?�6��&-?T�>w��>�f�?AL?Vi~>���<��=^Ĥ��T
?%�<�\ ?�nռS��>�t����N[�������?�͕�>���3]M>n^�������򂾨!c�6�B���-��.徂W�>��0�<�׾�?�p�"=��8�)��=�">ֹ����=h�����=.��7��O��	=�oI�<����ܶ=��a=���=ISD>��=�'== >��^>x(I�H�ƽ@��=�T�nۧ�����Gg%��	���	W��#���3�Y���(\����>h�_0�5�F<jm>mp���#���ƽOL>'�>{9$>�XI>��>��I� ��=b����R��]��<��&>�Bp=����=�}>�I�=����!�
�@�����;�ml�Ѯ��e�r}���ђ�I��7>�E>���=v����=��y>��'>�O��J:=�ԩ=3=D�r>�x'>~�>O�>�,>]d潴�S�]g�=D�)=�Bý�W	�E)�=��q>���<d�h<!�=�1�;b6�K���.M�U �=�o�I=i=:�>�7��(>�W7���>�i�>�<�>�}�>D��>�+��%�%���H��=V�C�o�}�cr:�ۛ(��x"�h��6����*=������)���Ǿ�=��G�>&[|>���>�|�>u�>��������=%>[=F��!��~�=�&N>lV�V�"=���=��>�_=��>~>j�\��K&�z۝<m�=R����I�<���< �<q>[=�����>�
>�}��e�#�'���m�΍��=�v%>~5��
W<Ry.>�@">�+��k��=H���v�=TM�<��&��1O�=����Q���n�5��=�	��A���߻o�)>md>��˽����1C���ō=�̽��=�J>ފ�<�"���=��=��|�3��_2>H��=ׄL>`����C��SV ���U�����Q�64���2T�ޱԾT��<U��=�&��M2�>T=��>��<J,��ۇ�F5�<+%V<;��?!�>&>�g&>{��=a�F>BV���<�G��j>��l=��_�X�?�D>ߧ��d&>��H�S�:}��<${�<��>|��=3eA��0m;�M�>�R���ս�
�/H�>C�>Y~�=J�`����>��>�a>Ϧ=��>�<��������<2��>�?S�7�i���<q�a>$)@>����,=;-ӷ>{J�8u�>_h�>nW�>�Ê�ϟ�>��>��>�O�,�B>PC>�n>0��2ƽ�����|޽�p����Ҿ|�������u���)�p�{��<�ǐ�q=�T�=�!�<e�R���<�U��e&B�0��<� 5>0>�_��V�=3X�<�|;�Z;���;G��=a��
�����5�E9���ʱ�r精$㋽Ϗ
>��6>S�U>����=�->Y�=�eV�4݃�Ϙ8>}�>v�P�YG`���:7���2=��z=ld�=���>��
�M�N���k:Pz@>�WƼrSX����C��=�>^{J>I�~<�/W>�S=�� >�Ώ>�h�>���7��\<�I�;(�׽�bv�������=�{�����ߓ�0nW�őo=9�=b>��S>��b=��O����p��=c*�r�`��Xa�k�p=�O>��_>=�� >�����V�pڡ��cH�p7>}bG��i�<��=XN��+�N;�@�]J��t[>,0�>4W?>�xp>�#<w���U��B9�y�=N*��?m�<z�c=u�f�Zo;0N��Y��=�+�>Ѽ�>���>��>�@>Y��=s;��/J{>��=�8D�����<V�+��ӽ�?���R=zC�>�W>̾>��>�y>LB>R!˼�}�=G;�=�ݟ�%�N��3�;+c3���=ii��V�yq��|(�VЄ��s��c���JCJ�y⳾2��-.���A�������� �=6��<�"��WՉ����ɝ彈+��Y���+�"=%m=����諒k��:�ж��+��� =��G��~&��n�=��ɾ9J���]a�X����I����<<0����������=��<&p��ճ=�0)�1:���G���D��/����5�Cp��.G�>"��<;=��>��>�)��;���
�<ne>P���4���м�=*
�>�V>뾽=�m~>:�Q>'m�<�u��
(= �>���l,1��$���>(/˽O��b_�,�+>�(>�N�=:�!>:�:�k�˽U}���� >�C=�>�ɦ=^q>[M�:b�<��ܼ�TS>~_�>��M>0oN>��>�ʩ=��M>��
>;��<\>���=V,��2�s�ѳK=`���~
�T��7��w�ݾr����¾���-�=>���W�j��<��=��%�!B���i4=�}ּ_s�;���얞��g"�OIֽ����Ͻ� ��|a����*�C?,���$�R=
w����!�ѵ���2{=w�-�� �=��>]>W�]>�#����_Tf�E�u��֑=�ק���^�.l��e����b�=�J=R-��)�d��X�[�v<6m�"�#=�*+=�v>�>it��I���@���Q>�Ƃ�j���߽���`>g\�=��]>���<��~>����<^��寮�A�M'2���M���<(Y���	I=M[s=@��<����N�ʯ��~ L�ː.>�j�>J,>fd>NLX>��D>�&>�>7�=!�}=K��=�P>�7��h�����,���jƼ0p�<��C�S9���H>+���4��!���ỽ���;I�=��������*��<4 ����7\�>? Z>�ɡ>悚>P�>�S�>	��>}	1>���>˗�>�g�>Jp�>wP�>�f�>cJ�>})^>��/��o=�9�>���>���^zq=>�L>-fL>otf����=�e->)>
�{�ذ��5��oZ=�~���᾽ �0�2��� �2�!{F���3>�﮽z��;Y�=+�=�Q���w!�����Y�Q�z��=�u!=k�0��9�s�<2�>�� �܅��o�-=�6�;�=��<Rz���/{<_½�����)�z�z<;�н�)=�&��ð��}M�<
��3о��!�H����>�>5�T>M�N>�����݁���=�A��L��<ּ=��.=ڂ���=x�=�mB>R#I�;_��G���"%˼j!c�V�_����!O�&C��(����W��yݬ=)6�#�뽒>/g�=9����V���=�j��]t8��k�=_G>��H>��B�&�	>�P[>�u>�c��Fx�=�j =0kS>���=>3A.�@��I�>:�I;ݶE>*��=�X;�L޷=C¼�>{Ԍ���)�����,Y=Ǻ�7;���{<�N='�v@�=�Y�=y�#>��G��&=�}X>H�"<mf���;(n>���=�d�����o���?Ͻ����8g=F��=NuX>��˗�<3�J>��;<`��D =�B#>�ɒ<�v���01����u��A�<�@��A=DR��#<����F>��=���=0�=��*�K$�=x�>�^G>��>���>we=x�7��濽s)��.�<��=��(=<Y�=eQս���������t;H,9>��q>�N*>��W>*�0>�m'>�>lӃ��X>si=�@�=������q=��=>���=5`@�3�ڽW"O�G]�����rB��@.꽕�$�E
��r��h�=
��=� =o�n=�>Η%>sv�= #���� �����iƴ��T-�:kj��7-�̱#��o&='���������;!��<=;'<D���{>�զ>�׍>v6t>+!>�mG=W=MI%=G�E>L�ܽj_�F�f�-��=畁;S&���%��2>�y���=���;�ܬy;M�����=E�c�f�潜��YY!=3���"�M�%�<M������M�����y6�����^|�Q ��F1���Z����<M�i=��~=�y��-=�u3>)i>�?i=6Jc��1�S�c;v<�T�ھ�|z�g#�����m�`�{'����Μ�~�ھ���8�����<�'辴�)=r��<��W�|z�>{,*>���=��>���=��2��A<���̉>��'��p���v>5�R�5�ۼ_[��o#���=���y��zɾqy
�0	����f���Gr�=d|��k�����1]�>����;\�ɽU8$�.�X?V��1��ڜ�Pt񿌾�?#�1?���>��H>{�>��Ͽ���y #��X�?ݑ?��@>s�=��$?���>��h?MF �5fڼ�]ƻ�r?�"?�\>Ĕ1����>�g�����W=S�d� 6����ʿ�ҹ>��ܽ���?��F�$<�?g��L}}>ܤA�tM?��>)]{>-��>�ws?G>+�%?�$��,�Z>t��l���*�5�`�о��G�-w�?��x�zn4=��9?[��>�$�>X�>����ֽ��P�(sǿp� >!o�?О���m�?xb��-F?�Õ�A��>9�~�O�>9FO�'�w�[]3��'�Yл��+;>�L���`=�;�]����=�)q�@Yx����/>�u�8����&�MQ?:�3����>w�j�1�q���=�8�>-���wO?B�2;�&�D%O���S�b?��5?z�?k�>NF��&�+1h>ݚ���ӿ�{:?�Oƿέ�`��^�h�޾�J>l����<�>�;濼{��2�澯7��"��=\����$��@���C�Ǡ�?�r�?��=��������Rkj��B:��X���?��8��?BY`������~?��>�i{?�c@ �F�7f9���>M䩿]��?�G�=O��?��\?Q������?-8��K�>�wq���=�s
�L���f׾��t��M�?�;j�֜��#r�>��u1�>�ۀ�{��?l]Ӿ_��d��?����'�>�x�?��� ���U~�b^E�URp?�K�?�n>��?��h?!����!�ڨֿ�4���2����>�^��Վ�=!?>.�>��=�IK?��s?G�?C\�٥���^n�j�vſ�̍?�Pz?t�?�?�����]��1�?9 <?��>ѿ(a==�~��L��>(�I?���=_?�U?>�Kn�j��������>�ti>ˏ��Jt�?��;#-�>���=��i�/�&�X�8���O�mW�?������>.,i�OK�?'t6>(���=�E?���?kxt���_�B��o�Y?�0B���?��?��>�#?=�$����X!���N�7"�=��ݾ�xy?)�i?\��o�7<7?��˾C��\���;�ſ��b�'?LH+?� � ����=�`>ԍ�l���k��Ο��6�D���`?�r��0���>q.�?��҇�>"�&>[1u=�˿�p�>�Q�=�6?�]���=&@
?��>w�Ǿ6������׾�oG?7_���A?��e�=����{?�}D?<t�>j�$>��-?T���Q@>��<�6?�V�?D|�>�!�?��?#�p���=}��v/#?z��>��>��d?d�ƿ�ģ><�z�5�M�N����;QY���`'>�蘾JX>�<c��'��Ⱦ�萿I�k����>�˟?Yn�?��?B2�?��q�%g��L�=�i�?y���0��= a���?�7_>8�n;Pw7�8��>��F?|l��Rȿ�>X��-)�pA�����=�N���^�>�a���>�;�^=H,?XX�>J>�?��?IL"�>f?�����B?e�U?�t?�A�?�wU��N#?qD�?�/=$�/g?��h>�@?���a�?t⚿�L&�� ��K�>,�?Y�W>�a��%�?����9�R��6\�=c$����̦y�����������1>��?�$��7¾��?�a��/[�e�/g�?=R�>��*?��>�׷>������?Z@⟂?u@�}ם<V�>S��?��>�g��5��>+〿�8��~n��\����c�4��޿mǌ���ǿu�"?\����dj��t<��n�v�>;�]�eZ?3�!���>O�o��.�?7P?+�/?"�!?����M��:�=h*?� ��>�N?��>���>��(� �{?|����SD$<Xy>�@�����?Q*0?�U5���ھ}>H?�N�>����%\ݽ
����g5�A��|�۾N֧=�}'�k)>��V�-�>��L�c�{>�ϩ���*�������>.d���j��=Ff(?o����m����T��>$}��2�Q�-�=(<�>>�����m�n�����?���=��V��&?=�!�1@~?)�/�7I�:�	�6���FA���x�>��ۿ���������m>�:#�c��o�>��=�Z�?{]~?�?���?Py�>0�>P6���%&��Oi?҉L>Ұv���㾣>显���*�F�:@��?^'�?�Ō>�F?���>���>�́?�O
�k.>t���پ��M?9�?I�K?o!��ѿ�˾?�����{�Wn�>��`?��x�=��?�����C1?��h>��n?E^�?<{�?Y��?�S >'�W���>cfK��¾�u?N���>�z8?ȝ8?EG�n���n�O����N-?�E��_����7��Z�D� J�?�X%�yײ>섓�B�@id����n?��>�"@��M��� >�/�>���?s�>��U���ս��?g��r�&?+%M?�v۾�J��(
�4R?�l�?&uI��u쾱�H>�ϱ�Yc�)��?~
�>��?7c>��g���������$>\��>zn<�@;7֌���ϓ|���D�<g<?SZ�>�0�?���>[(����?����?t��Ϯ�>��5�04�����=������n�>���>PY�>.7��.�?j�>��>�P'?\E?�l�>�{?[i����>��=1M�>7�O=]~Ͽ�"�?�]?�������<o�?���>ܓL>!�gH�=��W�����߾i�ý��������н�kٻ�0��ɾQY?Ac�>�?�]=�?Da�>1��?��=�n�>j	?��V>qn��?��f�?��@S�f�^%�>������RA?pJO�$�>���>�8���+=ƌ�>a>�v�=u�,������������>&`r?��>؞�?�V^>E!ǻΦ�?�n?>Y��>�_�?(�-?t�?��>L�;?([�?�7�EP����>�V'���4�=������$9>\s�m�����<�Hy�7q���?�l�?��?S�?�%>�2��k�?�ﾳ%V� 'U���A?Y e�6�?{!�>��>2�0���Ŀ#L'@���<?�\㿿w�?�?�ސ�hZ׿֝?&Z�?4�j=�G�tuX�'8;?!�A?68��-��7.�������>"�[�N�>�'$?]�?0OS�mn�?ш�Z�,?&A��*?��>�/?*:Q�^~=�%��?��>���?�gz��?�_Y�CYܾ]�?s�?�xN���_�	�ʾc�\>�v;����T>�J�����Ԩ3��4?g��>���HE�����>�
?�BR>�t?��7�=�վ�%�?Ͱ��Pb?Z� ���N?��ľ�W7�R孾�q��pb=��|<��ڽ�É��<��K?e�K��e���\#���Y>z��?�6=���HY���q?�>� f?��>�(�s��߾'=��`�?0dU��Ջ?Nh�>��?b9��� ?zFK��$�>_���V�o?��$>y�[?���>�ۼ�|���Ǔ�Ř��Օ�Ne�?Q@>�P�=��?�������>��Y?��+��>�	>o���ı?W���?�"�>�?�m`�8�М>�����>k��>�2?"��?/G?���?���ƥ�(�1��<�T<�K�����Ѿ��(��+�>�(4�`���K�?�޿�_i�ȹ�>�F�v�?�T;��ž (1�T��=$��?t�6��N�?�'忡|?���<��I�#����T;J:
?���=W�?��<�x��l)�&"�>�|^><ԛ?n	����?ޔ��5֙?C��>��>����B�>��>g⛿�ܧ?����+?���<iR�>$��D;�?��	��)���>C�Q?���{�W?1(�?f���>(���>Be?y�?hC���A��ُ���i>7��>ua�z��>�=���=�ϥ=�v=�~d?f������>+>!y!���?m��ݻ=��?!+�?H���q�
�~�>���?�%�K	���Ծ�Q?6 '��-W=���|WT����ɮS�Q�[?���?Y����?,��je ?�W�?�/�>�N�>��?��>�H�ےL?�0�?HD�?k!�>f�;?*��?���>������0v�P��>=t?&w?�D�Ҟ�g;��9�>D٫��F��e��Ւ�>֦1��f�>�*�=m�?�l"?��T���/>Y�5�F`?���>w�8?��?�w.?S�3��?z�p=�褾����>&�����K�?U��<� �H �>�~���i���w=��>z+��@=�cc�H&S�О��f!�7�?���?9����h?��>�T0?�����᱾�a>�_j����.ź=�L���>=��������>՜��;��M5��Zs��������>p�����c�|5�L��� �ݫ���꿺Q�<ߝ>�i�>��>���?�Ǿ��u?R�p�4-�>O??kN;?Ȓ?݌���%�;�0���o>�	�>R��F���u蔿C���'���*Dm��^\��n;�. ��'�����>a}L>a�C?�e�>j�>2��h5��J�N?�
�?�e�>;I>p�>D�>�Ϳ����?/@��r��>M�Z?U�
@���>oy�8�a?�νP&�?E&�?�=G?���?G���gP���6����?n~�?+��= ���S�%=�w�>��oo��?F�>��?7��H�?5.��U:>9k >�bX�nP���w>^>ؚ>�������>�?���!����G?C�?Q>���ɷ?��￉������f3��B�?~"?@��^=r��>��ܲo��O��yt��1?\o��s?Z<>>29�5;>}�=|<⺛;��?�}e?c�,�8��*F�j��W�
?xy?&�m�s�?ֆ�?��¾I�����Q�u�'?o^�?��?��@�YG?��ܿ#�����¿�'�*��A�ʾOX?^-?4N*??F<Ĭ�>����V���U0��p�?�I������+�]�@>Ȍ��2}?A	#?��?�6�Y�A?�!j���[?��=���K*?���=�'�5��?_�,�����g(뿴�U��M�%��p/�>�$?MQ#>��6>s?�"�/?:��?K�P?�-��8o6?��?=A)>9�)�!��>F)e?\�]?��B���=i�>�>��쾀��=�ҾNSľ���=R'?Dn�>�#$�/�׾�x����>��m�g��_��{=B(�=�
�?�{>&S�?el=���>��?�<��2��a��?��Ƚ�~"��⡾iy־��4�P垼w�=xJǾ����q?@,�?Ų7?�
Ⱦ�b�?��?�`��y>���?��8>��>&�>��?�P8?m�=J��9z�ÿ�?W;��&bi�4}�iַ>/Y������,���V�z�ɾq�><��=��e?���>wdI?1��?a�? ɒ��w�����b��9�
o��ߞM�tf޽���Ã6>��b�t�n=g�T��b�?pX��(]>N��\�f��e�>qQ&<ȇb�nڌ��@����&�l��>���4i@>b!�=6�e?���3|?p ����?���>������=>J\0?>��=.T��""?�3&?����Dya?i�?�t?_���S�?��'�{?��'���h?)�H>N�>��H�����J.�3�>A�>B9�>�E�>�ގ=}2
�ԥG�_�>i�%�S����־��]�p�1Q\�* ��9����?�/?UI�?>��?ޙ�?o�ؿ4>P��9�?�?N��?�7j?���������=.i���N��S!?M��=.��@୾��d��v>WV����q�Ù8?!i����5��?�
�? ݆��p�>���=C_y>B�?�M�5�.�_�q��T?.�?���?�=}��>�s���:������?nv�Յ�=�"c��7���xؿ��I��;�>n8���@?I��=�%���?�"�?( �'M���	�?������>N�K>�����a+�?�ξ�%��呿�~Z����2�Ͽ϶ʿ�4����; 6���Ք�tְ���'=奷>x������s�>�Ӯ;3��
_Y��z<�ȿKu���̽�3?u'�>���=��/9཮3��L5�|<��㿋ן��1�
`r��Ց��=�=�?�>U[2>���s�,?����P ���>��>�� 3>���>�����A�?��0>|�?�5)�_�ν��a?�@�?��>��?��m���Ԝ����5�?�E�?���?-?5��>j�?:}W?�|�=�Q?�^�?�ɾ얋=B=>�<���>x����>l�^��_�?�V�=SR��0Yۿ�n>��S>Y��?�'q?��x?��>�j��$\�>�y]="�>����F���;LK��3��>$��yT��ڸ�=s���4H/��s����2?�-��]뾡�Ͼ�*j��)o���>"s�>�⍿;�O�ξ-W�?�����>�j�>��8?�u����>	�>��M?�x%�-4��EVg?L�?tat�v~=5ph>�x>�z(�A:)?�D����?����W�E�Z����;����f�?�ϽL�?O��#������=W�q��oJ�c-L?�?�6)>�]�ޢ��4��I!ݾ�SU?i��?��?����m?�i�>�,�s+����>O8{?��Q??B?�u����=�������D�?.2?u?+G>Lz�?X��? �?�+9?��+?��>?��?�)?��?N��>�4?{�?�ד�Y����?�'!?���*�>�^�>������E��>W_�>���>�<ſAR�=V���a���_\����=`k�>�����l >�!�?��_?ec�=[H>	?CQ?'>{�� �">\��=)����Q���	L?<)�~�Ť�^Ĥ?4�b�6��>î��|���VW>�z���i����?�cP��Գ>�*�>�{�b��*���i�>5�>���-{>wn��?s���?������k?,�A?M�4ƹ>����9?�6?s�S>y��?��W�~b}�\�>��>|����h��i>x�����'wV���r��I]?`��?�P?���>Z�D?��?E��>rC1����?ݕ��h�j�i��=5�#=L�齓Ԧ���F? �˿��?6�o?��?[���S�??�g�?�o#?�濑�Z��>�9C�����r>ZJ�?��h��9
D���G�b�m?hC?䢔��J�?�F>�ֽmL�>�F�?〾��־P`�?��6����=�A,��?wy�?�xc?���lCr?�=�?L ?e�>m?^�3����>��>2l�>,�->s��>d�}=�}=�!j�?�@���>�V�C��?y$?��;���^?,֑��q�?hY?B{%>�"���	?�?��8��ft>��
?��ʾ�ȃ<�;#�F&i��g|?x�>��t?���Rp]?C?!q?���B�>�� >�|�>.�¿�\��:�=��y��B�?���?�������"���e�z��?���?wߴ=@�?��>��w?��5����?��>��%=�m�׌�?�#?�Md?�q���Z�>V�����H���V�!>sv[�rb�>m{�=/��?�%�?�b@�9?iߎ���=%~?� ?���VA ?a�H�ĵ�N'I�� �>R	z?C0�=xD?�I뾢om?���?o#=���ݿ�IW>B�0����C�E>[��>���=9�=�
1?���?�ʸ?PAj������b����ڿÉ?B��>�/��׃��T�$?#{G��,H�?����o�\��>"��}��=�yX?ݎ�� ?�\��JM?F]�?��?�;�����X��ۆܿ�B��6?徸������Yk>i�s>`��>�l�>��� ��>!��>Z^ݾgT?����RZ?��.>P��<ƶ��+ӾXr>L�$���"���?�u�b�?�m<�9�Y=�I�������J��k�����?a[A>�]�>Gԅ?paD>�?!@0?��o�A���Կi>R?f���J�?T��>q�>sq��
�G�c>I�F������ O>;�&�Ģ��|p��� T?�#��y����)��r�?Ҽ�?T4?CQ�=r�A�@��=5I =���;�����@������<n�z>D��:݂>xѽ40��_���x���;�����>dv?к$?��?1mP?dq
?���>�D��'{]�^��<�a�=!���E�ӽ⧰��������I�<ʍ���i��op���6���'�m)�>r��=��>�sM>��> �>�j>?U�>�X�>m�>
R�=� �~]����96>nV羰��>�ǯ�gk�>k�6>�HѼvM{����
��]�������(��^ry�����%���W'�xN��$-O�����~$ ����=��>-;�����>�f>0�>�� >M7s=�q>��}>[�D=s���9��π	=�㽾;��G���沰��	I����O<�%�=6��=�h|>Hg=��Y`ҾF큼br�z�>��>���=ިX>{�>��?=?+7�>���>M�¾$�+��Ƽ�!?W�ݾ:����=S�=��Ҿ�I�=q���"&��{��eݾZ��^<I����1<jL�������澺�Ǿ�vֽ�ơ��E��=2�gó�AK-���ྼK���|��{��=�
C��r�>'
(>*�I�We?���,_6>� �>|W?6X�=�Ca>^ =�<�<7ռ(�$<2P�><�O�p-��`�	>����^�/>��<Gᚾ�ν��U=����z�>�ѳr����>[Fj=]󧽷�н@�x��$>8�n�p4�=��D=��Q�q�=Q�0>gj�>9>Z6=�D>ck��	�>=O1��=�8�;��i��_>�X/=u>�>=�7���ϼ䕾M�#>�-����S�A�N�'T��4�=6F��q��?�B�d5�=F��KUn>T�T=��>�2>�8�>���>��>Ґ?<�(�w�꾰��<KD����>}-^>42�>T�>V��>9�m�֣w>O�=��g>���=�*�w/>f+N>�?�O>P�=�uh=�=�3 >H#�>�7��0��N����U^>�D�}gӽ�:;VC�>v��><O~>��<>ِ0�V^b>���>,?���>��J>��>;�>G8?�:=�*>���>P5h>�W;>�>�]���?E^���N����>l�=?m:�~��=�=@���|?=�?�m&�>���>�&�=�����5��������%߼7Zy��t����ٽ�*�}�<P5̽.�;�~>��>�g9�vD�>w�>|;>��>��=�>.L��g�>9H$>�$�>5ԼY5L>��N;��M=n�	�oa����Ѿ{��K���t�<����KN>Ql���d>��ݽ��>i;ɾ<o>�>Q��K�>��>&����۾S,��_a�=x��>=�=�彩pb��J���K>���9���<��K��X>�O�=}[[>n�=][�>4�?%�?Z>2?a�>��>A1�>�?A�>��r>ڔU>�>~e=�LѾܱd�0�}<_���J��2�Ӿ�C>��;��1���;<�JT����S>+}5���'>8��r:���E�y�>�/!?ο7��/�=�t�>x�?2�=5�i>J3Ⱦ*��{h>/�[����=��?%�C?@��>�?T6?¢ܾb>�j�>�/V?������>�.���i���>9ӭ�Wu=>C��>�0�>Pr�>���>D�=�D��׎=k���o�=�C�#�F�*��=Om =�eB���.=T.�>tT�=Q�>�Y1>�L����>#��=R�>��?���>ǥ�>!�o>�%���4���ڽ�0�H�]�<΋=��>�|>����9La��M���KȾ7f��������rSB�$��>�2�<-�z���u���o>3DŽ
�?�̠����<y�=<�s=uM>[��>ke�>[5�>�Y�<�`J���!�B�~��eV�_�w��Y��&�n�j!�> �<W��>l�p=�P?�E�<���>��aN	�%��!4��M����=K�ܽ�d���ӽV���<�Q�j��a�[�,�Ͼ6�ƾ۰�ó��wu�a���z!�K�W<�zF���=q;*�ۀz=�9��E��1�?���i`¾Z>�����L@���ݪ�]|���8��7��=�0����V�=߫;��v���Û�!쥽���[@���I>��L���-�������>o�$>$�4���Q�D>�=;#�Z:�]	���þgm.�Q^����#�M�����a�vW�L
�=9]�;�L�P��,�Ӿ�_����>1l�>�x>d�7>�V?�@>��?�?��t?�<��C?w����m��N>� ;oE�>ޗѾk��	}m�Y�ྩoJ����/	�F����W=��ݽ��6�>>�=��=�Q�>�G�>G>�]^�$x�u8�<Z�~�F���%�؆
���F��7���_ν3��W����>=鬾:Q+�j&��=�=��=<� �.#���������q�eE�49��R䇾�߃>Q�<#���3L=z����=1��>r�Ra�>c�/�s?�ٶ<��>F&�C�=�I�纊<+u�=��Ҿ)��=&T�>,�x>}��>�
�>^M>̴>�^%>��m>��=	�����>0��>�X?��ٽ��j=֦��D�����>!0L=t��;�>�<�>R!?��@>�N4��v =���=Ɇ�=C�W=��G�\s��F��<�\@�0��>=5D>��H>b��=w�>���>�à=B^�=� ?��>�?8�5>�&�>w�?�L�>��S>�n��`R>�W=a�u�Mx��|S?�!w=�sp>P�q����>�d=��C�3���ެi�����$��.d=�P���C,���I�������	>yuj>�g�;�5�=�>�d�<�ͽ;=�=D{^���8�cח�^_>K*E=G�>!2�>�'�e��>�W���ʝ���#�i�,>wb[�Q2�>�#@>�F����0>��F����>5ۛ��u�=~+�>k|>�#�>H >��=B��>/4�=pK�p���?_;=Cq�>�r?s 1>�j��E���^:��G>��8�呸>��O��Z{>ŁL>S}��[�k >��\���f�V��"��&��e���Tb�[>EO>�b�=��|>HKg>�5=&j��E��<�G-��:D��	���x�M��>�c&���<˟h�|�?QEN>�͙>By���">0�d>Q�C>����bC�8�Y>z�_>��7=�->ո��eA�U��>!1j�]�S>��>�Ѹ>o��/�>�0
���=c��/޽�9�=��%����>��=ȇ�>)۾��>!?�=!�>y:!��>?J���=^�u�u����޼��;x������֪����=d ���V�uH��Sĩ�Ҝ��$��%ҽ\�~>���=bJ��t?�������Ͼ�PP>,4F�[=4�	)�=Mʼ�gɾ>TY�Ů<>�] �M��u���e=���>����^�F�	?>sR>3H�Խ�=�!r<�o`<�B�>�Ƭ>�q�>�V�>w'n>z$�=I�>	��>��>h��>�>u �=��>�B=��^>��5??:���d<���<gｽ#=���]:�=��������?o�׋\����=|�� �v�6�F>��>W(>m�n=�>�CO>g�l>��=�w��
�>o&0=
�g>�\E?ֶ����=�?�}W?��O>�o?�cL=���Yt>3��N�=)S
?Nλ>��\>��a>"2R�K��`~n>�{+���4�ʴ��eXP��X�9��>0�=*��w=��.�M���.&�{'�琾~J�=�l`��!��Cվ^�j�����pz�=5���������N�'��+��3O�s6(�hV��e>��>�>ãr��6�>��O>CU�oE�=tc�>��=���>BZ��O����y�>��ܽ��>daܾ�蝽��澜 A����s���"�<�vh��/���>R笽,6ܾH�-��/&>�[��/>�6�>�Z�>f�>� ?k�y>�In��'->�'�=�\�>3�>������l>^4k>j�>��>��7���Q��r�M�yb��t���@��De��N�nƾК>c����T�yR�� ?���='T=>�y;�~>-�L�5��*�?�j�>f3
��j�i��>���o�!?�# >KE�?�^��u��?�� ���"?�2t<}K,>%�>�k]��2U�x�ɻ>鐓����?��1�Sm?�)?�@q��L�3O���t���8>�YB���?�R�?�p�9ˠ��)k?��=Ź�����; ��o����҆?�U?�s�=��?��=��#?;�O�e�>��B�0?��-Ҿ	�R?�_������]��~l�<�C3>�S�>?�=[�B�����{_>�77?W�>�1?w߉?ML����k[Ӿ�͝?�6A?0dW���;����KHU���J?����m�>J��?/�?;D3��H���	�>RrA?�Dn>{۽��>|�����1������So?M�߾;s�_�?kH�>��>Ʋ!?=�Ӿ
 �������p��>L��Ʉ?>��?�ת?˲@��*�jq���+?x>*�.������9�e�?$�=;_��B�>,D����a���S�����>��Ҿj�=������Jl�?#ed?���?L�>��!���F��F�>�h���6��i��:4��о��S܊����>���?���=uF`���G��b2�]�?H��;|�.?Ґ?�����c=��Ծ9��?��;W�@�X]�m�.>��?⶿��G>�oC���ʾ�!�>�����@�>�K">�������Ň
<���>AJJ?Kʱ?)��>/֗���>�)C?���>��(?p�D>-�����-R?5+,�~u�>�+�>���?o���ֺ���U��p[�b�^����������@?�l_>��>���>wS¿ӛ��X��)�E�˧?�䉿>%��J����>"d�D?A���΀��w�?��T��`����
>h2��N*5=�al�$���=�����%a`����� Ur?�
�>6�2�L��>�2����>;|���;�-o?��?��?xvp�3�۾���?yrR?3�*��#�ry�?�.G?Ik�>ZV�>vt>φ(?�z�L����t���O@9B�?;�� x;>l3b?����^8���?C�?��Y>y���>w�>/?��J?��??Y�G
?���B���:��?Ő8��>�������f�>j ^���6>�D��#?"e���L>c��*Ɲ�@j�k𰾦ʽ���?���>�ž���?���
".>� 6�eb�������?uF5���ѽ��<?W� ?
�?�C�<�V�U�=�~Ͼ���6V#��u��'O?�J�<뀏��G�I������z���a۾�6�X�?�HX��2`�e�~�� ��#▾�PR�y]4�1H�?�З?&_�=lv���(��5�F?�ZԼ]�P���r?'�:?aF��2O���?��p>A�?�'�0��|�>.p�=�>:4���r��X�?���=L��>ax��p�>�Ͼ.��� .5�QB/�[	,?�����s�=Ί�>���E)=eɗ�� 	����*K�>/)ξzmu=c��?X�2�@ZV�WF}?W���2˿���>��?Ɯ�>���LA?���%ɔ��?$?j� ?Z�?�F�?��1?o���3FQ?��;?��>�쩿���>��>��L?}X�?m���I�?��t��v#�4�;\��=q��>AM?"g?mvp>�O��D��F�Ǩ�>�nL��]�<�!��B'>����=���>]]>��j��=��L��l�=��>�)��Z��>9} ?�vϾ7�>j�B=u���C3>�'�>��Ǿ�T�'?�-@?yo?XBI?�Q ?�(?�?�=���	Q��v�����FX��-�$�}�>�*	?�C�>����A�UQ�02>Q~u�.>�~(�!TȾ�@48L�*ǋ>u�>�!��>}Fþ��d��=�p����;�!�.b�>�X�?��_@��1@:�������("��E��(F�>�}��2W��מ����z���?`L?�>��3@���E�&6�X�X?� ���e�h[)��+�4�_?��徛�	?�XG?�{?9�~A���^>B�s?����=s�He��B%Z?o�;���Ͼ�bT�؞*>�h=-�>Wf�>�Z�>���>�U��u����>�ߣ>rH�=p�	��?���>��>	��>k���P�>���=R�����r��yO?�y�>δ]���L�(?�@��� ?�ܠ>�9"?��>�&�?���=?����s����d7�>�ބ���>I��?ΞM�ᰂ>@N�?�� @W
���n��gb�>m"s�`۾3c��m�= ��' �L�ؾH!?#.�����1?��=�����Z?�\&@��"?Ǌ3@p�N�Q8�>ϻ�>�as�5gO�+~?����I+п�ؿ��:�j����>�]�=B�*?o�T?i����>#�B<�# ���[�Xz�>|[*�gi*�Q#Ǿu�>4ʱ�J�i?�O�>Ǔ�>���>��~<�=�����c�?�S	?�J�<�.�v�?���>�}?�
�>^Z�=�+>r�������ҭ��ͦ?j/:�����,?$B�>[[��Ǌ�>"�C��M�Bp�<x��s	?���?�7���Ҿ�I�0��@�<j)�nVI?&���i">�b�������?w	f>I������>���>|��?g+���m��ꩿ�ں>/j�?E���ľ�L�����o���b�J=&?�'�?2�?5[�>�6¾��r���?�/y�*����>u�꾷*?�5 =FC�?Vp���}@>��>0�"?N9������I>�8>��7?�^D?�|�M��Z�=��.>�؇�^�7�G���=O7w>��A?��?��?wƾUп=>��ֶ�>��;�`�>T�4�^�ƫ>��>��>;Bk��9?E[�=U?����> ��>�q?�gP>8�Ǿ��?8�J�x�ֽN�����?gI?���?=:��Z����> ;��?���p̋?���?��?��o>$ɧ�>��>(AC?0ˋ=��A�s�����>x�}�c�ɿn0z��:�?�#�?�"N?�^�?fF?Y%?ߝ�=�w�;�mc�.��<��>sm྆*̿a��?*u�?g@澸��&G4����ȏ#��ӽv(=O	��sVD��?�(�>��g=z�?�{D>���>	/�=���>�M�?xk�>M*<?�h�?�[ �^�F��-P��M?���RQ����>cEk?�������	��>DpO=&1T��5�>�(u?�x3?r(��D{��>����>8��>�ux��mc���R���>�⯽����殹?$bF�kC>�����Ҵ?����Cϻ���?h~��;���+�2�>]�?�`L�Ҩ@�?FI�}���/Y8=hv>�Q�>C��>��F?�w�>尒�}��>b�����R�߽�>��>]y?62���wV?g�׾ģݽb�<��t?_�B?�}�>ȣ>R/���:���ꤾ��JI?�7
�|s?�8�>�s�?y�B�1��s4��B?C��>�4/��TO���>�[��U�n>������?�v�=���P_@�f��>k?���?�O{?��b�^V!?��@	fV�1����?�r9R>���gݾ��?P�?b�?ƿ?�!a��Q��NP@�5L��w>�K?���>q���e�6����>��S0(>b��Zܽ�����,-?Ɇ>�6�� �=�븽�}ƾ������>���>0�B?UΛ��>?sFX>����|-¿dw�(|?�?!�?N�?�ݿ??����
H<�R�U�:zh�!s�>� ?��,�
�>� 
�S�*?ُ�?��'?�'?��?Y��?��?o�?�d�����l=�-G���>L�?��?E�?��ھ@[���pl�^$�bՃ�v�d�T��$�G?�r�_��0L_?�k>��Ҿ��>6�>�|?���>��?x���F�>�>�#�{�Ⱦ8[B?�7d?%�/���H?v��>�o�?o��>m�~�1���<���>�睾�;Zi����Q��q?��>*�Q>hL?���F��>;���>�\��}�������dѾXL�>�,&?����>���?�u���xq>�
�˹b?������a>i�>K�/���=������
?B?�($>��c����������nӿ@T�>H�2?�
�%F!>�:�>'��?����*I?*l �w��>fΧ?�ݬ?Ul�F��$�>2E�=`��s�>�Ќ��)м��>H�=�	?���>_��*�����辻Z/��'?o�ܾ�7�Cɍ>Z�پ��>0����O�����?}ز�m�پ�2�=wq1?`�S>t�<@�?�M�:#ʎ>�_��AN��|? y1�>P�?0�K��}
?�}�>���?�gs>�kD�q.����ż
w���"ؽ�?�=R�����>�R�?�0�>FIe?o��� ��Sg���q�l!+��%�<a⾜��?LS3?�
��Y��=�f?��7=�>@��c��&�� ��,w�<]�F��j3<K���GU�>q1?�$w?ch?tt?���<���/�>��>?Rm?򁣿�H<���J�:?�?�[�?8�U?�I~?!NG?�j�	[X�MT���?��ݪ��%6���'>�,>���,򾟟7?ќ�>_@?��C����;{��>g\���@��U*;M�����;�]��Y�������b[�W�i<�����Ľ
�߾ܲr���R�EE���Q��>�����{�77�t4�*�=a��=9>�m��R7�s��)ξ�Zz��~@?���=1Y��+�>�X ��0m?QY?#�w>o�(�����`�>�(4?�,ɼ/�>h��|�)Od��+����?���?��=��>���Lc��Z%�ҕ�>;�K?r�����*>uv�<�!�?��= 6���=C2b=��=yN��P��?m��>�F�q76?�ڔ>�Q��1=�d����9�m"I��U>H�+>��$>��׾��-�n�Y3��H}	��3��qD�>���>�B��)�~���}?@���$�>.�>+E�>�c�?�z?�iܼ�����y>���� =?�P�?�`?� ?�c'>P��>Т��L"?�X����"����=\(�?���iﾙF,=��?����3J��߇�Q�&?�#�?F�?eO�>F?c?�ʿ?�O�?�{?��A?;�Z�����K��"l?2��?��?�E�>��e?��}���>�撿|�}?[�Q>�%�>�c�>u�`>�y�>l�X?Z���ac?6I��y��?��4�?�Ƽ�|��/?.����E�ٮ@?�����V��_�=��?�Tg?ۘ?B�?h�D��`?��Ι�/�Ҿ=Iվ	�q?�}���:?f���q�>CO�?�0?o��������η��)>gJ?c,B>I����/?����Spr>v�?bEȾ�_�x��!,e>|;	>Z�>߯b����?��>�$.?<� �D{�?ư޿q�[?s�����ؾʫw>5���XjR?($t?�󯾹-���IY����>4 ?m���B~w�xD?u�[?OS�>eNF��P�?���DE?ֵ��hX?R���	� �D����\�>��־�?p�?^��d�G��\������z�>C�M?��>P��>�}6?e�0��L����o�Լ�>�=�eq�C]�懥>X>$
!��Џ>;��><�?]� ?�Ĥ�P���{�==�c����?�G?�� ���?�q{�4D�� ���thW>Hi;�؃?��>C���1�`>����}�vH�>V�H>ۢ������o�c?�̀��Э��l=��!?/9:��&�?�@��Ѽ�V�>2�=�d�Ȕ9>�����1>jtվ ��TĽ���=���?vVI?憙��K?����r��X�������8?c��>���>��p�h<9��a?�� ?_�+>^�>�$�+u>)�}<b���0�>4G7?����ikK��?�?��k��y���w6=�ӛ>�UH?�/i>�@�J�Q>�Q�?Ʊ�=��e>?�;^ZJ?�?4��>f��=@?[��?r��;�>���\>N@}�����-��rvi�>�4����Z���:h??��6?�B?�e���K��\v�\O`>J���ʊ�>��>�A@<�#�=�3v��>�9`>;ِ���>wH���io���Խ�����򗽮!�<؊�<�s?�V=K?��U?��?I�~>D_���G>�4�>�C=Y����'��Ӄ���2>X��8���HCk>�T�>�
�z&���?o|�>3���̶�>*���e�Ŀ�`�?-�J��"\�G�>�n�����ۄ����ԍ>)��>¾��ݾ>�E?>���>1�?n{B�Dk=Z�y?g��?I��>Qs�=d¬?h����*����������o�?[�� S������{_�I'�>����W��?��>cH�L��g��?���?�j���.'?φ$?���>�۾�Ħ=a�h��~���"�=��>�(M�M0��0�>�f�>?�I��x"?6�><_
?"��>������=�I�vش��Tc=� �?c`���=�ĕ���?��<����=cT;?i�?^a�>�U���"ٿ*�>��F?�|\�� >����%?����8��M�?u{�>��!?�&u�m�t?�9޾*��)�!?�ݭ�RP�=x�=~�>����qfB��~/?�{}���>']���>�;�ios��[>��?�oy��
=���>-��>�	�=�4Z?1��>E���q�<o{j���A��M��%a�/◿uF��� ����>D�Y�be�>�b�=_�?z������I�>��;7O�<
Z�n$ ��;??/k�p�r��a}?�>?:f��p?��[?��?q#�?`N�>eX�����>U��>3?3?%)h=ɀ>�P>}��ի?V]�����=���>��<O��b����0�j�1?$Ty;���侢W&?���E�8�M��������>%�d����=~�B?�^�?��?\˄>L��>{B^>L�;���=#a?.�&�U�;*�?kی=xWd>Q੾�����!�?3@�>��m;9��>��	?��?�O�?��#?b<5?�Қ�w�?+�ɼm5?�"/��i��12�<|½!�ݿ��~��� �N ���3?[��?�H#?F�5?�;�?<J� �����\?��ƾa�O?ct�=e�?8���o«�J2���>Ѩ���4K�F>�f�>��wl�>C8Q>?���O@��?�����?�U?��T�yO��;wf>-������i�Z=�����)�ov?�25?�%@��<��V�?��z>�S�?Z+�$C�?2��<��5�wOĿ��#@ZQ˾���F=���	A>�q>k��?�����T���>#2��5�?*�d��c�>q�����1�/ #>��˾}Iľ���q=0��>�3�kP?sd>`о�`�ﾫ�2?��վ`�sls=�)�>]4?��+����>$郾���y4V?c�(�#Ӿ?\w&?'B�>7yڿ��>0�h?rm�L��>/�i?s�?�'z�G:=��q<�ڪ���">İ���$�0웻A��~�1?��}?�ϣ��׎�j��p5�����|?�{���.�?;� ?K�>ݢ ?��0=�?O	�>�X�ң��h`� :B�_P@�<�����>��;�∽�S��9=�=Q�Q?�|"�1�>��?b��?=�ʾ�봾�q?�C�����ŧͿ4
�Ś���枿��?;��JJ����>�C>6������>"->7��f>�>�Q�<8�2>9�J��wL��žʿ���v� G���X��59>H
��&ؿ�ȁ��@���I>�[?B�1=�o?|?Ogr?9!�=??�~�>Q�?��L�<����3��;��ǐl?*U��?�?�P\?):>+Ju�I
?D�v���������=H�#��fR=W�~�2���I�?s?��.W�����6W
�
2辝�G��վ!�!�7�u��E�>S�4?�y�?��}����IeJ?��>��>�`�>5�0?��k�|��ΏO>�+�>Y�C�X >�S8��.R?!��?Pc�=|M���[?���=�����Y��t�J?h`e>��[�6����7?9`>��p���_�s�辘5�:?�?�f�SS)?��[�(?Z���<�?��K>y0+��-����t涾�0��b�>h+����7?�����Ġ>g a>�T8?79���4�?F�?,��=q:?=ρ��M�4�о������T�3������>Z��=�� ��A�/��=�*2�+�6���s?���>a��>��?6�S>Z?��>�??1�s?��U>QN�M�>�@,>n>��"��ʉ�+�>�hf�~'��?� t?Z��������p���>>��>@��}B��>�>F/?���=-���I?�QR��?>�?9�����>�H�?�=�=����g���{4;%s���;�e˿��٥;�����:��H7����o¿w5�4!��>	���I�>���X��>Ҿ���?t�#�<g??�a)>�h?8�>4P�>��j>��Q?y�>Q����5��v�>�BU>c��A^�� 2�h�?_�=�mϾ]�I���l��p�>v/;��<>������6�h�q����>�U>�D�o�`�E�?o�-?g�1?�t�?u���F�pަ�� H����������	��i��<�G���j�r ���P�g�;�vI�εP���-=s�?�X�>���>�r?��G��S�(��=�XI�!���T轶�U�h"?~�c��Zy>cP���e�΍>"��>�Ȫ���ݾ���)> �⾧p�>��1>E��>k�i��h���`=`�ƽ��u=��s?�Ϝ�`�ú�>'�5��B6>�N?�¤>�?K>4�>�>t�K?�W��]�-?b�־l4?�4�<iNf�$�̾ 9C�(˂�M�����k�^�����[�>u�8=#��?�*c�f2)������=�>>��=��z?|C�>�(��?�(>0G>np��S��}���X�=�'�=�[N���=��
�J�Y�N�>Rc><i����V���=�>�Y�>���>��=��S?>Kw�=�f�>�RE?�2 ?Fu�����>�:>pE?Ɍ?��>qs���o��$�P�x>��K�u�>B�b��?��n=Gm>%�:�@]^������>��)?G@��@���n��)?YD����2�b���?r��>���>,,��ܕ?Z��J�2?�r=O?�2
?�Q$�A��<�)�`��>h0˿���քB=����=��\�>v�j?�1��'w>WJ�=�g?����b>4��;�0S?)V"��� ?���>���=%X���� �wξ�˾Z	q��}[��F���1��h���q��齾��=������>��	���?3��>�a@?c�?�w�>���>Z�?V�?Ch���"���c�> ��>����x��\]ݾ:�S�FW	� �� u����=�R����S=�-�>����^ �?��F�����'z?e��>��x�Ί�>�g?)gv>z�C���2�'�����>�&>���f6B��	V>)�þ�'����,�ɉ^=�Ù�]Q��C�]���>��>��!>����?��?[��>�1?�w7?U}���*��� ?��>{X+>���*�w�<@���}z>�����y�O�7?h�q��=�	>�u$��E�������[u(=�^�=�ƕ�)�>���=�a�a ۽�g�����>�4C��8C>|�>;�ý����n�>J1��le?�ٽ���<��f?�!?x��>�G|?�%�1;=k�a�$"��*��>`Ι��8��{�>�g�>�t?�L�=�$�>ޟ�=���>�`�X�V>��>6��2N���9>����=ξ\�5�ķƽ�	o=��.�HbL�l�{>�U>G`?B�>?�j�<.j!�N?�wG>f����>L����R?�>4?��?�)�l�X�%#��_=�|>����R�5��`��u@��BV����`�,0#�5��Un���M���i=��1�b�,U�b�M�A��>�(=\��>�Ƚ��V?23P��s�>��5?��!?���>A�־O��DH���6�>����G�<��=.�g�I��I�>p�E�!��>��3>C�]>\�?
?���}�>/鉽m�y�ׯ.=Z��
����u�#
����>�k��tq�,R	?��{���B�J�e������+��[پ�;����s�Z;?O4�>�d(�ÀȾK��QE�Z[x�y�:�u�����8���~�M���>�x��E��Mx��*?,>>Y9缻���T?���qm�Ԗ���=�E ����I�L>N-j<8��>DC3?���o]�>����ⰾf�o>Ky/?4X+=��>%��"�'>ˑ�>C?U6 ?��i��[����s?�m���/����>���h&?��,?���?bu�>?�}?��.>i"?��?�+?�)?�қ>Rp?�Ա?�h>�ҽ�c�?��Io�>�#�`̘<]K�>{�ܾ%0h������!��(�\>`��>Ӻ���>.T?�"E?���?:B�ci��W������4ǾF0:��^��7���f�R)�e��=�s��6񬾳P�>��*���S��>�P���8�2�/?	0>�ȍ��½��>ų��|l��7꾗�?U��=0��>宋��?kK�F�?E%��OLd?�T���
?��?��0?�,+���>��H��ێ����i��<?�Ѽ���R8?���>�q?�[D=���>�.�?H�C?1�v??`�^�t��HH��rd>��������þ����&���2?7�v��K��n�>W(,?�-V?�'���e�� ��6v?lH; >���;���K<[{;@�T?��>��L?O�>��V?��?;[K?66F?�Y?��X?S�?��2?��?�� ?��?��e?+n>��A>���$�#?��`��;<e�?Fne?J���`?g�p��m��(���=1�P��!������H���(�؎>�M3���<yu>E�>�̐l��ʣ=X�}?|�>O�1��d����>X�{��>1w=���>��i?Uu8?d��=j ?���K����g>H��>�?%�x>�·>�uo��e��8þ^a=G�z�[�Ͼ:3��殺���/�b�b�>(:�=ؕ0;PJ��s�?�>�B?�M�^Ď�mU?��]�U>��;�?�Ő?/`y�	)�C?/����>���?�%�!�X�d�]�t$��qD9�����c=	<�!�/�vt�=,��>��+?!ʠ���S?�����>)�ĺN����~R�e?�?���%�����=��K���j?�ܾ�\?dm>EL�?�� ���e���W�"�L>*@�E�n> �þǐ&���>`�?E����Oe�G�f�M��>�%0�+H.=G �>@3�>�Ծ�e<�&[8> M��,��W�T?U�o�6?6h˾�Q�?����=�.?F�#?�;>��>���4O���	���=�ι�ؾ��.�>���`>?ɓ#��ܼ��>���=!C����e>/�?���J���,��g���,���?tK�=�?�[�X�>/�3?�Q=>��">LX�>4�̾������??<�	?��0>Fq=%RI?�;?����w��/7?눾ǌ�=�+���i>|�$���?R�>�ҽ�/[?�<�>�f�!��>��
�t�w?n�>.m��j�Y?tn�?�@?&����r6>V��8�?�����L"��p�H/>1&�{�����>���=n�'=��?P?�0r?�b?�P?:��>w�?�+?2�ɾ
L'>'[?ONO?(w_��|t�@<���yU=������=��R7�>��g��SW?7�>;K���:�?=��>�Lh>U�?�b?��4?��?A�h?S��<��[��樽9N3><�>P,���(������>̀�=p�>�h�=3+�7��>�ύ�4P�=��X���B��3�?��k�F�H>��=���>-">�a7���>��,�O�7��<d��A
?�u>�x?=oM�>"�>I?�5�> ��>z��>R'?t�=.p�o�>�����C?5	�I0�=
��=�X�>Ψg�)�j?�i�>O��=�l$�t�K�[N>��P? 쾐�~�߷J>�����9?�]-?���?�i?�ռ>S�ؾ�]ͽ*�?Y�=C�̾�H(?1,W��.	?�7 >�l�T\�<Ş!<Կ(������t�h/M?��ݾ\�6�N5��<�=���}b�<N��FV?R�>�B�>��>�%۾㤿��:?Z,���ٜ��>�{J�G�����>��ɾ��N>�K��]�>0Ҟ��L�Hp����8?a|J>p
?'�9�e�����=�z�>F5�T�/?�w>�>>ox!=A9>�,�=Ձ켿v��(>I"���u��2>�H�>��=�L1?�=�>��¾`�F�5�=���P?A�N? �>C�? �J?�ۦ=�xt�n�?���=�+�=:@B���=�7�>�?�щ>��%?�������Ev$��@�=���àK��D(��P�1��)ؒ�o�>��>*�2�$�T��2?�e���۳>W׾ȡ߽��)=�e?�U�>ɟJ>�0�>��4>��v=���`~���?'�y>���<H)�H�\>���>�cO��M���,?�aܽ"�>8�=��x>A ?��=�W?fi}>�ȯ>��I��<��[׿��?ΧU?��?q=7?�"��MJ��]俁Q�>�����1��6����)`D���l��s��`Y���P�w6��i�=�(�>��+?>%j?V�A=��:?�߹��aE>u�?Q�����������똾�	�?h���N�پ��罢u#?�F�`�ֿ-�{?a}�Ć���U�=��ӽp��"�??,>E*C����Vy>?		q>�+>t���H��?m���P?���Gg�>Bx�����=N��>Z�;?2�.�'>T��B*f=A�=�5����2@����=�=�+;��;�=���=�߀?�U>m	 �fP���jɾ
䗾@�?s�7���Ͼ5��:b�W=������ܾ�Xﾄ�?j=��CI�Й簽�/�>q����~p����f��J��ܑ ?f��H|�>��.���?�됾s��?X��3�E>�H�>� $��>%-�F�`>) /��6?���?[�?|n�?�[A?���>eS�������S�>��b?��������J���<?��L>��m>�F*�g���C?S�{
�?�dS=���4>�h?E�.?�U)���?��?��J>�@?>��a�� �?���?���>���>�FJ?u2����I?c��zI?c�>:$y��-L>�2�>`VJ>��T�/�>H�J?)�?�wR?-��>US?ę���b쾢vh>�݈?Z>C�>�Ź>Zjl=��M�ED?*��?�Q�X2��g?E���n���C�qS�`M�>lT>�^��R%�,���V��Qݾ�(����J�uy�>:�;�5$��z?q��>�K�=�B��d��ߓ�p�2>���> NW;�jk>��˾���Pݣ����ŝ����?ԓ?T�4<��>{P=�/1>��.?�J�?g�[�����>��>[-��V�>�$%?@��?�L�E޷=�{g�|�r>O��eی���]G�=��)>�r!����n��>4hM=�V���[����%?�j?��_?.��>I?���4`�=�2���e�g�>pÆ�rփ���˽>$�>�w����>t>�>n�`�L��5���o7>���r��A���1'ս�A��OB������oK�(���?]	[?d�?B�$���6>��>+���i>ثP�}E?,?8��>�<�xϚ��=�-�?Vr?��?6A=C-��W�==l���X>ƿ�>��>�RҾ">��=�^���!��i�&#3?|��>�:U>X�?;���4g�6�5�`
�>YPX>�jR�X!2�J�r���w���`�����>/�>�?��>�}p?�*y=#�=> �?�$���4��
��8���4�J���-�	
�=&𾶗j?^�*���"�1�2=-fT�V$I�SVk>f[U>+�]>�����>N(�>�bͽ(�	��>�N�{��>��F����<ͣe����?�,?��O?��X�$ȾC]>E!p���Ǿ5�ƽ�SC?��?,�Q?�ew���&�~�	�N�U�)i�>;�ŽI����>KʽY,�>��G���i�����\E>��?_��?���=�a<B����V��Z4?M�Ҿk7%�����z�>;�;>���\/�>d�>Xa7��c<���.�ӻ>�(>��<Pg�>uk�>�A��³Ҿ$���h?���>���h=h׌>���_�u����C?�>�!=+�`>(��=�2�>|C�OP�=#�>$3A�Q��>e�>�	��ݱ�=	��(?^�?m�$?�?�%1?z�]?���=D�>� ��uݾ��g��#
�PCM�r���6�x=������>�'�'A+�@�Z��$V���|�@o�#��,@�	�>s�1<��<?E��>f�F�ҏ˾���>���9fu���=��>� .?d����O>�Ծ��+�F?|̖=�P*=�r�>_!?��B��3>'	��8��n�>��Ҽ��5>ae�ld�>�¾����WU�>"��/D>?�?y�>>��?!���v��u*���pw��2��G�gZ��[?�GK��5�?�3̾�ݽ_z�l_?'/>]#�Cw�>��?�ψ=
pg>�r>�r�?�>9k?&涽Ѡ�>��@����#'>��u?�M��0�>��	?K��>p���˿���žg
�>�1�?2�?�|F?��7��bھ���>U�<��>wn�>�<?e��>nÂ���#�vR��U	q=ǚ���>?6?+��(���;��=��>���װ���%>���>���?�x��=��#�����?R��*?ǍT?�y�?�h�?dǵ?��f>x��?�`�?�yI?\�?_Su?v2�>���>��?F�,?֎�>3����>b�.?:?��S���p�>s�?3{�Ӥ�<[�>�>sb�
a�2?9=bEξ�c��C�=Ll��2>X���t;��;��%�=?ɢ>�?����ק�����3+R��Ik��pn?�� ?�T=���?���=w>��?lh>�7T��ii?�:x�Y��>p��k���o�>��?S����c/��5�\m�>��	?ϱz�>
>wow���G��_�CK�8�"�D�?��>�U�>�9??& 4<jq�>q�>�諭�p�;�0?D}������b�=M�	>��?wB(��˾.��Dh��%�}�G?�t����?�v�[��>F"?�>��>��Ќ>�v�>0�(>�d"�m��>L�0=�c?��b��ҡ�O��=��?�־�Y߿��?4r�>)��>#���S���>�G?��;��!���?>�a>�->fW��5?�>��Q�ͽ�ޤ�S�־��>�/�=:D=*��;�_H=����I�`yO�����,&)>�>ϾЙ��� ����ھ�q">˞��1��7	������z?8u�UZ�
��>ڟ?��=��)�>wd���r�=M��W�1�mY��}ξ�Dо��� ���5?ju�h�+�aݾL����(��'>y��h>{�)>���>���D��=��>e�/?U�>B��>�S?���=���뛣����>��!�$蚽eH?,{��.�>�5�>��%?�[�?�=�>´�<O©?�2>9�>~fI?c﷽+� >��k?h�>����n�>�_�>=���ZE�QQ5?@$�=�X?j;�<��'�>��x#��*��>��h>M_?,���;�>E�)?L��ʣ���4?��J>WGJ?;���>�)�>70��>��G��]����,��>��>�Œ�dz�\w�>�>ƥ>�4>����s^?RL>���>�B1?Rbi?7�?��k?$i!?v�>eF�aZ���{d�x?&Z��"u�^/�:9H�=�Z<y_ھʔ"�!=�_D�?�k��V!)�����X�>�Ċ�@���� �	����>`����/��(V>Lc�����-��>m_(���>,�=���
�>xJ)>�C�>%CԾV��>:=?�q~=�S���P�����=2��qd��K������qI���<����񀦾��>^��������yp?2�m�F�7������=?ܭ�>�<>��X�۟�>gF�>o>�V���?��?�	��$�s.?��\>��D>4i��-��?Ä2��C3���-��������=b��>$���1�A��c꽂�ž�i��N���Ň�\wj��巽j�
�����͑��mL?�gz?�M?Gq��]h��UA��,��]�?��?��e�>	���`�?&�]�����Q�?O�>����{���'��$��"��/1��f׵��K�Y�C�� 3�,1D>b�?2ת>�S��:\��u0�&����?s��>˚
?��>ӭ#�Zr��p:>>��zӽ>=�>��?�:��S��>�F�>#c���B\>7�@?	/>�×��>�3��K��ǣ�K�V��m��eH�>���3=�`��'�>{�M?0��z?���>χe��Y��?4��=Dg�?�q �� �DǕ�[�M�_X�3,?��#?�މ����?B�T�;�㙾��r�L��>��L>`U? �=��Q�Ot��ې���?�� �:�+�>Ai�=��>��L��()>��w���?�H��O�=k2?
[��>u�nO!>�f�W[�Ջ���I��?���>�'?J�q�\��.ޙ>	z?@(¿�Ⱦ��^����1G:>���?e�׾i�#�����{<���?�y�=΃�? ?>h�c��2	پQ��=�|<>��׸`?pȐ=�_�>�lP?Z1�>tξ�O�>7u��|���=C?��:�Ľ(��=�T4>(վW��?>OǼ'9��ٍ�h\�>8Xо0U��%�>xHU���Y?� O�iz?����Y�>3c�>�o>������q�Q���h?)��>�����c�>Yu?^���4�7����=iҰ���>Ĝ���m�Yl��%����=��_?�*ܾ +�>�"��5�>C�Ծ�!e>UQ�>rּ?Ra�>g`>fA���(�<#���\j޽m�H����>�����t?sDϽa��&�C�a����z��O�?ҝ>y!3?i��>Q̰��?�B��H?Ǐ ���>|MS?/r�?J��>�C?�M��ɂ��k�>�s��B�S����>b=.?�(���"ƽ���<%���KK?v���E�?	��F��?2@��	6?�%򽱈�?�P�Ch>Dp6��"���n�>w9�>���>Y&�>��>V�><r��X_?����ݙ>e����i[?'z�=P���0{����>�nվ�u�>����m�<�:V��2S���w&��D�į�t��=TN�i>�Y�>Ĺx<�ߍ�:;?+�����>��Ѕ�>��ھB�����3����>�j�>T$:�Qo���-?���K� ?�@�?�k?�6�?�o,?b�?�jT=̒p?jh�>�.?��r��Ss�G\��-��=5V���q�>��>�:ԾN���s9���>��9�{R ?n<�g?�랾u۫�1���X���b����>��=��m���.�K��� ?�$�>]7Z?W�����>"2���g?����d�>C*ξn?�+�2�%?)뾑@?��3�C>;��?���?mM�?�w?��A�0���Կ'����O�|?�'0�Dsl?�!>uC�x���Fq��Fs���5?�8W�c�p? jU?��R���Z��Q>����/�ǻO��f�f>�r�>ѣ>?�؊�-
�>��o�Q0�?�B����>�*��y���b�`k�?�\-?D̴>;^�>��r>��??>� H�XN�>��@?�6ؽ���d#J?꼑���I���;1�����>�Ċ�l��>�lؾ�j?Cf�>SDA?9!@>�o%?���>~�����>U��=̚>�T>�u>ޯ����J�s���U�����?5!v?�{�?�
v>OZ4�	k��#�q\�ae�?�	�>��|<-v7�����"�C�l0���tp>꛾>��>f�'�E$D>8��w��>�4w>��ȿJ�u�R�g?}� >�Spb=�@��ap?�z?�>�=?TC� 娾w���Q9��ſ�[���M>B���_��>�b>4+8?t?q㾹�޿�i����o��da��`?�Ծ����;Gۿ.�2?6��?�~�>���p��x�վ�<��_�?QF�h�IR>�_��@$�>B�=fU�>]����[(>�}�Fk�>p����\>����ʢ>rཟ�?X�K>G�#>�vd?Ii�>�TY?�����?8�$?�X=���R�	>���=�tN?���>�&?O��?�g�?���?�V`?O��?w��"��j�>n�w�p9=?�	:��K�>����O�>y�>U-C�+�=�Dl�p�>=��<�o>�>����&���Ҿo9�Mֹ>t�,�?Y��ڞ�>��s�0�ľŅ�>��$�d}��ٷx�e�?���?)9~?�{��'~����>��=*���#����Q��(�˿��Q?0�"?17R?��R?l�L�vw<���ߤ?��ѽH� ��W��.��)o?�=8^�?b4�?���>
M?�r�>�ڀ?��ÿ_P���F�8�4��?>�Ow�LWH��?7�;z��>�T��h��>�\�=��%>��?�56?��B?�=��@��?Uz��i"?n� ��*�>0�I?�a	?=^M�
��>le�=C7q�mO=?+-?�#���`��忿�%<?vDR���>��>T���%�?�$5��b-��X�?U�ɾ� ?�]u?�����u�>ÒB��T_?��7]2�c
�=򸧽�J�<��G?��=?�cU>�SN�����Q�˾�� ��Q�>y9>7�>���v��E?+��-��Bfg��?�mF>��u��?�N�==2d>7s0=>�g�����-��v�����JA�I�/>�)�=�d?��͗���L��i<ܾ��%>ïƾ҃�>(Q��=呾҅���@?��t<���<�4m�y/�=�|/��7��x{?bv�>�?����#6�?���=
Î?ݵ�>U�E>��?��gs?���>0��?Pfs?�&�>�+'?���?�#??�=��?���>W��=:'k=�#�=���:þe<���M�?�k>�y�Q���?�i򾘥?>V>,~�=5	p�e��O>�1?��]��kg?�֓?�B��)MH>��F��M�I���i���$�]�?>��?�W,?EZ��f�6L���?�6�	9�?�'~��4�������?�h?Z�O�E��>�7�>�Ծ���C�'��ݜt����?@'�=﬚��&�>��>FM����7W��GȾ�w��]��j���J>�)v��X*�:��>��>��t���[��+?oE�>��>z�m�[������=b���坿���?���e?�\��U����=�d�='I�?�J,?�ڈ�r<�Z&�="$F?)`�ky9?�J�=�Qξ�`��Sm���>՝þ����:�U?�� ��"�O,?��8��ٽ�u�>	G$�;%�����!v�,W��"���T�q�%�:i�V��?+�Ⱦ��7=��K?��ݽ;�;1r�>7��>�4�>F*����*>������ѿ���p�;�wľ$x������?G>v���h?��>��%?
��Ђ?�w>V�5?{'�@ϐ?g�>9�\�g�ܾ3�?g�?g��>�u��??���0�����=W��>,�~?���.��đ?����WS?�h%�� ?͒�~�?9t���<�¥>�;�>\�q�ow=�2�����=�����?y���*��>��.�m���3J?��һ�_�>K�>�O?y̾����8>4��;&>&?%�Z��X3�D�S#��N+>>�?oB3>�1�=nz��e�>��>,��=7�?h�	?M�C�VxB�;�+���I����:�(�IƊ���f>w|�>Xg�?Q!L?`���-��5L�>����G>�U?G&�d�>y��?��=�^7O?�+��I->cq?a�˾�'����>�$ĽQl�u)��|�>'lL?%b���5w>��h=n��2
f?�7��T�FG�~����#�>����$�v��ޜ;��<՛f��ڟ�����L���վ6d�o�=+�'�s]������I?/�?Wp0�sSþ�!�>����>J��>�Z>k:�?�#�?P��?�w1?�Z>�?6�п�bE�ɤ>��z��J?�J�>��^?�2��O��>}�(?���h+4�P1�����?'*���-�=�ȫ>��>��ͽ���#��
�?z���]��y���c���ql>˛b=pʙ? �'?�����9�*��wɾ}����>̼L=�>�����Y��y�7������N^?Rzi?\;>?L�m?�7D?U�j�ފH> ��<�>�9J?�-?r��>����R��b���|�T��5�꘾!�>��]�dz�>E�c>}.?��+�ڵR��Y"?�*?̶�>�mI?,�!?��?ą�X«=�,�DϾ�e/?�f�������*�H?�� =�t��#�ݽt��>LZ�����H�>4H�˾a�;E�����7�1��[�>������d���	��?� �?��?'�H���?ʡ�>A��L��=���>�8ѻ_�	?<�>$2�����9>"1�=��F��c���^��:�>���<��U>�>���>qE��оj������F��=�$_>N@?��X�� Q�3Hľ	a�>�?�͔?ƃ}?cH�?n��!��vD?��ݼ ~>�)���>�Q������/���żZr������F±�`YܾӉ��h�?�%!>P��>��Ͻ��<�=�����$?G�>��F��Gp�|a=8���3;>I1�8D�>��&�X>�>�r�>�X�?��?-����ؾZ~p��M�����]�?�{j?�i|��L�p�R�!��5?3^��==�K5?eY�>�%��s>���=>��t��W�>>
��D��?��������	�v�N������#3�0˾��?R���j���l������ǵ>�=�>�V��%��:�ξ���X�ܾ�?�X^?a+�>�U���Ą?���lb��&)4��;?�$��6=׾򾸔׾![4�����F?���7�X���Md��E��P���v�>�@����>t�8>�S�>\FU?�f>?2?�)=:7y>P�����>F�@?0x����?�O?��;��D�>�ʟ=��?�5þ��1��2���?QK���ल>�N)>ϫ>�'�?�L�>@�$��P��/����Z?1L�Q�?�??�w?\��ċ>@1?:z?}(�>���>�D>��9?z��>$Q�=�ў?�t��Ϛ��s�վ�EX����>�@�]]=��?Q?:m�bm�?�?��U?Ě�c�m?�b����<��d���>s��?��=?�x��@�����>��>����w�ƾ�^B�kW��M��?aü�A������M��>#CU?�>�>KE@����>SÐ>ו+�ݏ�?�3?��?�"_��,�>r�¾���Y����A?"XZ?^�<p���(�u��$��p����Ⱦ�~2?��?$?Eż�a?H4D��HH��a�.G_>%o?�.?L��=����>8������>Ƶ��?C�>:�?�� =`��C⼆G�>r3��ZPD�P"�B>�?,=���=��>���>.[%?nZ+?A�_?S}�>O�R�0�]���?V�>�v&�� ̾_��;�<[�b�%���9��!����=�#���>�c>������LB���j�>�C	���վǫ^�3C1=�*<
X$>�1�>�!>���=@���)����9�~�Ƚ���=ַ6>T�6??߽�R�݉�_�>3�5?M2�>G?܎�>"�9�S���9|����HF�>Iy�;70�����;eھ5,�i����+��i�>X� ?�s&?�k^?��>󢺾7��K7��1�Ӿ\��>J��{�=�1cѾ��Sy'��>�u�>��v>:<�=䶖?��a?�
��"v��}��%ka�X�=P��� �~=a,��̀��R=P���}㘾�M˾K�,��i+�s����l �3���tOv��R �W6I��9���&?�Q,��R>���Fr]�*�����y�H|e��D�ƙz?t�?��N>ZKW?t�=CL��$�d�5>��?�/?4X��n��J)���bg��CF��>
?���?�8�>A<־�h�A���0t�>�l^���{>� ?F +?��?6�ʾ�	�����m	�-;�>>��>��þ��)>���>�t��lV�>�1����>����u�<�h��/��>��S>��p>;+�>�B�>�xJ��@��7Ż9�U=�e����>�01�F%�><�H=6��aP���{?	�>-�<��>5=��L�>��:�>t�5����>&�~=�9�>X
4�9�>HT>��?���>��B?�ׂ>(�>�&۽Ꞡ?> ?��>��>d��ټ ��	�d����b?�D+?��������ꐿ��h��V���?	����B�=����$^�<r�H?N��>���>t�!?WP�>(��JԾ���<n�`?��>������-���1�|$��<�¾)�w�uG=��(�JO??e�N>L;���]i�vc�'8�>�/�>�v=��r���$0��d��2>QQ�>��F������F�8?q0c>�bƾ&��z����~>���>�h���I>��ջ4��?�����ͬ�N� �Y��k�>��`�%��>���>�?&Qy���y=��e>jmY?7j׾n��>�R?�?˴I>C�X?u�O>j�=��[�0��3Ҁ?�)?�+\���d=�\�K
?�L�?�O?�g?FJj?��=JvS=	>�<wm>>�x�>��T?f�>	N��IK���m��P�*��?�w�>i�?�.(�<�(?�>+��<|�ؾ{�{?��=����K�	�,_�����!'���f�a?�=X O���x?�>t�]?���=��E?t��>,�f?��X?D�?6?/1?��?3�?�s�>��S�֝�=tH�?2�S?����?Zݧ����=�I޿�W>��9?u��>�Qm�Xt������Ⱦ9S��u�=
����d����>�/���=�>��.uE���O���Q?��p��6��=���iN��g_��	�?w�н�t��U�������>��>���阴=dH�=�����3�>�='GH?'~�>��@���`�mu�� �5� ��<v�/�n���>c'�>����@;�r��O>� o?-٢?���>i�?"Y>�m>��ܻ�Nw��s?�A����ݾ�B����#?�|�=u�g�'"���1>���[9U��IX�{}�䠟>�O�_-/��L)r?j:���	?A�?��L>�{6���þ%�j?�
K<��5��Pm���0��ƛ>)�>�%z�z��R���)�?�Sy>�d���f9?�C�>��=����2�> T�>z�<J@���.�>�J>�@�?�?Q%�=kѾQw��􇭾�þ^~>(�?I�뽇ً��T�5���X-����>�H�?Wٿ>�ή��6Q>a���������vh��l?1�?QB���w�L�Kn��2<�z��<���?��,?�[�Q�8?�ﱽ1�དq����>�6?0�W���&��?;���s���g��/�~F%�ED?d�[=H���=?Bm�c?���I�>��?ZE'�?��>� ���C���!�+$�� ��]m��7�>��>�[�?�~��A=���ѐ�=�9<Vޟ��"n>ة�>EOP=F�����?^3�?ׇ�>�^�>��ﾀ=�>��\>c˽f/�u,f?��>�����N���M>�*����6�������1?�Z��i�>j2<?�ɸ>�)�>�j=���<��8?-��?� I>��?\KG>��=�ĺ@��wA��˵�� U���2"!�3;���5*�-1v>z�ܽ�nc���>�
�T>�|?,?�?KYa?w�K?H�l>QJ�>W�:�Nζ�h��>%�����=Ě�>F�>��� ��n�H�Y?��.����+Y\���>^����p>�8ݽ��>ƪ��F/�>��*��U�p�K����>���<����͔�)E�o �����=I����-W����>|���T?z���U�F=
Lm���?��R�d�뽜d7=�*��T&<�}�����>��>'�߾�,��n����(a>�@	�^�վ����?>��>$sY��Y���e�>�N?HK�>M�??�K�>��Z?)2?�rK��ۋ>�2�>�� >�+=jU;�=���{?׌���{��*�>�p�>��L����.K��v�>�S�MrA>Τ=�D�k?C���e���BT����=��p>��q�V@�9�E�ܵ	�~�����^�褁=�x`�=�'?Y_h�WUE?Uj�6�>��۾]�>u|�>Q �>*;�>��ľ�A<�Y�H��3\>�b< W7��Oľ=&\?Wr�>ux_?҈�>��=Y�����=��}���=�j��>����)�>�5>?�M��@���z?�u�(��Cz��&Q?��۽��P�:��>�����?�[νVǿ@-W>�<=��WD@$ڐ��`B?�A`�mh��0���?R6���t�?X->��w?��j>#;���F���< �>�1f?��c��o��rm?=�E?&z*���"�w)ʿ�ym������>�e�>>�B�!(�9>�?���Tj9���E��U����>!�D��G ����ԯ�]��&��X�>I��#l4�K�>��\?:+?d�)?U����90?�5=>�7�>�E��(
��K�>�G��Y�C?�m?�9����>B���m�>DG��z��YF�pf>�����>y��>Fe�?�>�>�~Ҿ.�,�ȊX>�S�?���>�)6=Е??�ѫ=��E=g��>N�d=�+�xVX?��⾦�c>x�?p��%��>��m����?�R"����ڽ�a��#�?���;#�?��~�9�>�@Ͽ��?BXv�D��?I� �Q?�ҥ?���>�;�>�P�>���D�?������
�f��?(� ��o�=V2�>��p�ȣ4��۽��=Jg������n�=��?� �?w�Y?��@�̠��C�=������=3?9O,>/|��5�eE?���>��3�=
W�����/�Ͻ6�&>:X� &��.�4?��9?��1?B�T�y��?}O�I��>�r>4�?C�	>O��<3=�;�?��ɼ�G?�K�V��9�?�K��*�=���t?�@�>QO=zgN>Ǔ=zq�>�1/?^Rھᗿ'?<�l����*�>C�;�3�&�J.���>!����y�=	C.>\9�ڶh>����u�?�$I?�>r��<���?6}.?q��f��>_�?v�R?�	�R�����?/�M?��=fi=��c��
�����@�
�}>=?
V?�S�>Ie�HUt��'����/����?��@�?�Oe�\�?�p?&�!?!�
�E�?���>�p=��*��s\>�������j���~K�x��>56�>K��>�	�>�д��.��uU2?]�>s&��p2W���о�b������&&?n��>�x�2S>x{�9���J�Ӿr��>��R��s�>~.� ����_e>��?�c�>>x}?���W�#?;�>��I�bM?5|�?`_�>����b�?[�H?F��>~�Z?1��>D�Y>//�����?�����_G?c0����>X �>n�.?;���=惿����	sz>ȒھZv�nH?��?�c�(q�Lº>�l@j�@?"��?���?���ZJ��R�>D��?�"=�-2���&��x�t?}B-?�J<��氽t�����>�m>�t�?���
�z>�۾�	�	�?����6�T �?f�<ϭ��*>�g!��곾^&`��ȅ��;��x��.9��ܣ�?�A�Rw@Ъ�?]$��jK�?� ����H�V�M<���J��H�Ŀ��>45���Uھ�n�M`7�n�5�L��>�64�&Q���������"�>\a����>p��>����T�>��?H��?�gR�K4O�ѻ?��&�%����ܿ�X���Žj�>�à?���>~q�?_��֐4���OX4�΁���9=�@t]��u�߿�v�>{N4>�
@ �������/%�Q	$?[�?Ɖ0>��=�"�?�׮??�b�D��N]߾���>NN�$.��'���):?�֜?e��>Ζ@'�R?���?>��F�1��)�F@���;��ā�?_�>�+>|X���f���`��ʫ��?�����?�!��tND=�5��$q����z�!	�=�񺿺�3��?�T�wo�?w�[?Lʊ>����=t���W�:��I@>�CR�������½��=����x�8��ͥ�_���J̾�/�=�?J�����O�>��̼�_��ҕ��!��=��>��L��4�=�A6�{?j���{8l��p9?���?yҾ�]>��?.�/?u���,`?���?M䏿�F�?�*>\��>������B�нtGW>`g��C({�TT?4,	�CU�?r��?�H�?�� ��iL?�Jξ�cP���޾ť�?��?Z?���Pݿ��>�?�l��&�>��i?�~i?�%t��8">.�A?\昿Ѽ�?��j��u��KJ�	��9~��~��?�X?�`^?δ#�u��>v(���}>�D�?�R�>�y�?�Ip?�9�>p_@gO�?X:b�,�A>/p���j% ?X�_?ui#?#�l���*?�&�5"����.YG=B�=��m�`f{�@�+;��8��?HwY?,(Z<��8�vH[��'��B�?���<qɠ���\�W\�?��<KW�uxP>���?Sy=q2#?���>*�7?tF1�[fV?�ॽ���>�����>�k@���?�?�v�>�ч?�G��aR��j۾��9�X��>^�?Uо�?��s�X�>�|��k>?�yo,�����q�~�w��ڤ�> ֌���$?����C���:�	?�<B�yt?>������K�?�Մ=��)=�K�>�:P�Ʒ)�sTU�n�x?9�>Π��A�`>����r}���
��0�࿼:�>A��>���>�x-�����X�>87��N��V���(x��R?��4��/��Bz�?&:�>��?��a��@�?z=����?��>����?�P8>׮H>�lB��bT?�$����>cf@>2~{>�6�>��ž�?N(�?`��?,I?�s��a\?#"�?D��>iS���h?�/a>��K��&?�%ܣ?4��?�><��>����rA�?��=��)���>�%�?�z?뻗=�$?�3�޾�r<�\׿�3r�����ظ�bG���>h8�>��\>1�&�Vj�茿yT�ʽ%?rc��gp?F9$>��㿛i�>k�����S��+��� �2�����=au��P?{;�/@C���r?M��>� ���{<�I9?< ?�[>	�}����S�?��g�y�f�.sɾyЌ?w�'g��.Qt�<9?s��<~`�������?Q=�?
_$�#�u����?�jI� �(��#��Nz?��s�f��>
��q?S���д�j�i��w�M����9��FA�|�U>��u��q8?��&>Q?�kҽ��F@osҿg��5z��t�>p\k��u��;�K���>#�>yZ���| �P��?�a�������}>�w�>  �=x���X">|	�>^7��sȼ>#��?a�?�����?��Q���\?s:�>���?uD���޾o������#[N����>���;1�ŏ�?A�\�����&�D?�oV�r�0=\���o5�=�b�>،?�8��T�2�»w�N��K2������J~?�E����>Qo�>m�o��ؕ�X�$���d=��>*q�?�?�u��� �ݵ>J�$?�(�?X�����?�q?�d���l�<U�����=��.^5������5e����l6e��b�?'�=�"?�@PQ�>\� >&�T>�  >d4���X@=�.C?Ԝ�p피(%���?{Iο]�?O��=�0?�?�i����Ѿw����ah�̳f?/��>т���/��a�}��N2?(����Ǿ
�M>��W?�No?jSG��p��Eą�b|3��:��$?����>?���؈= ��%�%��4�?'�:=��>��>�` �Ol�=Ԧ=�^�>���Ӓ >g�?ZƊ�SL�>�a��O��]}?��U�N>�e�=%�>؞1<�p澚�?'�>?5�>��,>��t���s���>���>DE��{??����Ͽ<Ə;>��������������?�YֿQ~l>
�h���־]S?�9�=n���M�>c�]?����W=�2��u�?�?"��>f �ۮ��S?+ʹ'�_?���𡿴[v?�E���!?��?P�X>?����$��o�����?�uZ���}=(@	>B!9?�hK���;�g"�~H�?��?C�?R����r?Z_��B^���T?`�>�69?�1־K$Q��݊�aZ���=𸩿���>ڱ�V�R����=G�½?3������E���gLB?��?��*��풾���>�X>?X�>�,9?.�>�����.Y������9?Kƺ�:���#Q�>�L���M��/�(?�@+?�,�>9�	��Wǽ��S?Zb >�D??���ڄ�?�i?�Q?1�潂��>��D?7�?nV�ʤ�>�?�E�>őο������>� ��'*I?�4�٨��I����0�V>�;��� ��8����5@"<�<�V ��A����?���=*�d>�>��a*�?�?�
=?�����y�?�p�>IDi����!���}+�dj>�%6��圾�e
??2������o���O?wS	���c�Y�>�1>���?|#�)�ؾ���>M��>	���\O��/�>>����G?;�?�5>A��C�ξ2��?�邿�,̿��ƿ%>�?8�>8$g�9�X��*<?�"I��,�?Y���s~`?���>~�?�@?����0��>�-N?�$��I���H��>��a���>�$�?5Mp=wP�=	N���́�80�?�� ���?��O?�
>-ھǸX��j5?�4�=����R>��1> �����,�&Θ���@�?;��ن��Tv���>X>L�������˦��Q�%��?k�þ��L��3>(�����"߀?�L?�*�R�п��U��fz����2U�]V����2?���?���>�k�>X�;�j�(�WS��݉�y���A�?~���⒁?���=���>��о^;%?0۱��/�?z5?��]���]\�>�'<��> ƿ��^�j)վ��>4�>נ?~��%X� |=?E]@�2�>o�?���y��>�.���7>t����37?Q��>�$��6L?���>�mҽ��@�<?;����C@3ǿ|�_���������AI�7�?V�!�(ԅ�Х�?6*���c��ށ�tHm?�2?�f�
������?�9F?\Ȍ��E��`@a��>"��R9[?xE ?`w�2�R�(ز�!�*�̓�i�ֿ"���m>�_�>���>��}>��@�:T>�Ш���>?ξe�?�h>F5?4a[���h?�ܐ��D?�c��0��h>��>�h~�m����������>�<i��~(�g�q���?���>,���V>Y,@R��=X�`��V���n�=���>q�?�B���J�>�'�>�lG?�Q�>����V��o	?��;�>�?@;�>[��>i�'�d�U�-��!\e>�?Nmν0g=?R���\�t?���>�V��B���1?��v�?�*L��%\>��^?�ƿ��>�^?��?K?=�>�o�?��>�ɿ�W���v;>>�j?�%|>\Ӷ����?S\������+x�>���>#�9?d���W��������lA̿8r��\����^��j��3���x���2�����>�#<?$K??����ᓿ��?00�ky���<����?oL@��BO?����j�?�,?@��;ǧ?ρ�����w������w�?e�>/����?+yA��V?�j�A;:?��?��w?�ؾ���>&����h<i3|��\g�Ы"?�(V?�aξC��=�}���>�� M>no?����է>�O��B�:�>�yO?Ƀ�PV��o� >�S?�"�g����r��F�QcK?��e>�q��W?���<�^1?��?Z �>�[�?+�6��ґ���<�@�=N���Q�t�<H�?���������Z�̙�*�A>� ?43q���s�ZE?bE�?<��>���=��i��mg�JH�it�>&%?�Qz��u�e�j���_#?N�*?�N��օ?ɻ�=P�> t{���>�;3?^s�?�(�?��S��A�z��n�7��%��+�?t��>,��=B��?�o?^E��������>`�߾�-J>�]���2���d��ݾ�0>ޒ?Ჾ>!׶�B�S��I\>�t>���>w򺾗PJ?�h��ʾ�BĿ] �?X�G?���>�>n��/?M����Dp��ȼm!6�37�75=H�J>hC8?^L��8q��Z�Gx>�ɯ>��I�U�Z?ƣ?6�.?�=�n>�i]���8�	�����>���$����q0�ž}?71���:P?X�:?r��?u���>?�O��N�����?A�;?�m�?�t�>_�>�`>�c�m?�+=�����ѷ�M¤�K��N�O����=!q^���Ŀ���=��ڷ�>;�e4�? �-�ǽsɩ������^��?���A?�Ƌ>z|��ͫ�����c����W>x'<.I��Nn�K�H���*>T�=aU?T�?o������Z��뾲=rs���N?�l?}��������p,?���m�S?U�y?(8;>�2������<�P?�Σ��j;���H?��ʾ�������>m�J?�
�P��>r?[1�?��Y�2os����?���ʽʋ�?�A��39?��?)+
��_��k��->�T@�����"��$��.�S�!���>u�_?M��>4�j?T��>��K?K�����ʄ�<ĉ?ҕ�?����2�\#��i�]�B��>�ao?B��i��>2]�>ϕI?9y�nw���(�=A|b?�P��߿E�EW��'X}�on�=`����8�=;m$�=
?��k�J�z=�;?� �>��w>t�=��?�Q�>�d]�4
�>��$�oJ�>rվۤ���Jn?* 2��_�?қ)�?s6��1?�IG�)T�?*���?K��c��;Ǿ��ﾇ�5��f>R�.?�é>�5��!�P?���?­!?T�?�?�?���?Q�x>��>?AnT?�O?_�*>[�G��`?��T?v����^����?c3>���,�?��>�\ꂾ����]�?�҂���?��ۿL ?��澷+Ծ��k��,��S9�#0�?��S�������,T?���>+6?k��?�n3?0[U=�t@��?-$������>$�ǽ���Ѝr�fP@���l咿J�=�x�$���پ$nx�/.��E���@��O>��y>�n?< w���5�����@_����\>�]�?��_?8;�>L&�X���֮�!n��5|�?u1�o!����2>?��?�M��=J��K�����> ���zp�>����?�$�?������O���*>Rf=��f?��Ǿ��?9��� ���0~?�@�?7т��rl�̱�F�@@``�=)	 ��_�>�S�>��4��9d?�<�>�\����8���
?��=���>����ㄥ����O�=�#�O[�<=
�u�>����X{?,L�?�e��-�eʡ?!S�?�G��W���+4���>�Q�=^?�6�?�A[?\f�����A��0���GW?[�6��^��û>�|?�H��}�ڼ��|�<�5�2�m^$����>j�>.J���)Ͼ��Y�GL%��\�>�G�>��q���>U儿�r�?tڻ?w�,?z2�=�K�?��Y?�0=�u?>�&�?��>H��,唽�5 @M�?�'*� #�=���?�ް� 	��Td��G[�Y��>M�{�že_=M�d>�/����>%Qs?��J=9�_������=�5?L��?{�1�nף�5d?�ϳ�0.E<O����\��l���s6�����wB?��Q>��
��]?�\?�฿��:��a=Ww?<��?�N�?j��>d�޿щ�����?B�=��?s����?�q��]:��q��>��(?t�5���R?�S$?^+>$`q�x���S�I6�lD>?��?��>�傿��>�]?��;<�����v��/��>΁?dE��=����H�я����Q>o�X�j����þ�P���~~�����7����>*8���zͿb��>��?F@V�Ŀ@;�?|������?��A�]>��?�J���))��*z?7bk?��*����}�?V�˽�S���7=?������G?gW��Aƾ�꯽�¿��V?ب�?U�2>�ܫ������ü�J��K��w��=�*�>���V��b��<�h�?'u˾QE+?b˫���= �5�ߎ6���^>�8��:I���\�2���j>��=��=?-����;���?|���g�=K��>H��>5�>;�>b�;�q>���>Uϰ>���>�%�>¸>i�>6���]=?���о�"���=5�y�☣>e��>eE> ���e��>A�V�T8�F�B>簒>!̈>1��>׫�>���>���>V��<�=<��þƌ��e�n��.Y=ب��]�=(�E>�Э<���l�����U��<���D���V:)���A�Mzݽ�b��-�
>���>7_>չ��9g>�֑>��>~�ĽB*�<�@�����>s��>��A>N��<:/�>u=>��G�x]ѽ�L[���I>\����\�|���=�">-q�����=�^ =yĠ�m����v���J��H>Y�>�7]�h�.�*B���ڜ"��B>S��>i�>.u�>�@�>�IB�$:��yu���<�>`�����ߠ��c3?�Ύ��E>��Ⱦ={��R	F�8�־29���y��-	6>�8=��Q=i�O>�Rl=���e0����>�P�%����@���_�=�l=s�B�c󗼗)�=��>#��7&:=�c?�7,�=q�=��D>�]>Ĩ >��<>��=:U>��>5�D���>�Q�>g���d���؅�h���<�|>Bl�=�>�Z�ݺ	=�>�ݯ>�K�d)>w/�>��1����K@��G¾M�־�+޾LW#��=i�P����k:>'��=� ����(��Jy=�,��2	���֌>�~�=�;�=���<v:7N��㼣>�;%�(�>��>�-������C�p��+	��o���hÐ���K���������>��=�S��L|��N�����z>8f���\J��!�<�-�����(;�>�>�+>�>?l��Bڵ�\K =*��>������=�6��<e��>[�.�m>0+>���&_<�>T=y��>��y�=Ӧ<�AG�+�>�O�;d��G�����q>�;��K!I�:I�=���>�m��EA�=� L>�,�>�듾�B������m>��H�O�<\�Z�uL>_� >�ͺ�xG��@g>���<j}�>bGQ><�>�Yx�
��J������>cL�'�=&��>��?�煽I,ܽ��ӽ�R���X�A��r� �u��T
��,�>��?�C%>m饾��=>҄ܽ~d��/�V=M�<��>P1�<KP�p�>�*���H��%�b���u�ؾ(�>�F޽!�8��5W�)w��:68��ҾS7*�G}����>{�X>`1��La����=+��;XL�>�ǽ��=�|�>y?y
��R<��n�nR5�ã�_��;�+�����>"��=���<�)�8�>��=c�v��4��]|�>�_�=.|a=�Ul=��>�h򽗆�=@��>?��>�о2�Ľ*�	����>�_����=�p�TM]>�j���'�ϾЉ���rǶ�|��=���>�_�<��X��f@�E@�=؁��3`���*<�&>�dg>>�=�{�=��S>�Ӿ\0��;��)���`��d�<��I���x_�m�}�k̾@�(���<*��=�a7=dw=��Y>�㫾��4zx��2.�+���<��E����Os�)�~�ک>�Z�?>�A�>��f>A��>���>A@�ܙ��	�3�r4}>�+:=��h���1��>j�^���8�� y��6>T��>]��=#)�>��>-��>�V�<��6���A��,b�L	��@�.������7:�'��:�(��`LM��3����߾�65��`�㖪�����߾à�>���=l���������=�_\�[š<%�i��C�e�>���>�Vľ�x�>x�=_C�='Xl>S+��J���>Sc�>j�=S�>a'>�����n�<!*�J����rվyP6>��$>QF�<p�C>8@��
җ<Dl�=Q��=kF/=�{�>��;>��ͽŖ��J���z�2�����>3R����A�C�+>T�s>�xн6�3=�!����=�ٸ��<�ݵ=Z�>
�=~�>��>uC�>A�M�V�j�s�=ܪ�=.n���e�K����=p����Ĝ�O�S����>��>[�>%�!>]����q/��X��7�=�>ޮ2>�������=[(��6K�FV�<�>��>	�(>�>�l�>t�+>��t�of�����=��R���}���<P0�=>���:>q*T<{Dy� Y�F���/��f�N�<lD�>��>��3���>v�>r��=��">��нm�<7�����>қU��|S>�>�v�!ZS��ܽ'���꾆M.>�g��*�˾������ �^˸��Y���l<���=ׯO>�q�>m��>y!�Uʾ��׾1fʾV��>nM�>��n�9O���>��B�=�fJ���~����>�_�>k�־4鈾����Ȍ=�D�>D�{���=�3�Ď�>�k6>��]��G�����>���<<��8>-]�>Yϒ���>�h>��w<���P�;ݝ�<|�>��N�S�6=x�>��>>
�y��Q_�_q�����z��>��<���'>x�=>��/"�;j�?���>T�;>_��>��>���<L{K�[r4���#Q"��tR=���ӛ�=��p���K��5<["+>�ݾ�>��>����鍾HK�����^���������>����52>��=�0�? �:?v�p>c��>�ǋ>+�}>Yݣ>�0�>;A>��D?�{;?��>���	��>��>�都�vľ
|��.����>�}����=���>+t?�%_��bkx�%�W��$��
�D��I��tm;U�u���>V�<�v����ϫ>�#<����s�����Sbi��c���<>0��>C��>�!�;w>�3S>��)>Z|�=>�ӼPA�>Z�1>mnA>���i�W>���=�rd��@��=gN�L��k�L��LZ=�:�;�|���w�?f�=s��횾i}�=p>���<���>���>���>�~=�4��ԍ��T<����
mA>�Uu�n5>�5�>�R`=�BI��<�*��_���]n��'E�p�ԽH�ξ�վ��">2e=���rP�y�ɼz$�=�Շ=�t�Z��x��=F�=���D<��j��m'�>5N=��"���>	V�=��4>�پ�mb=Ȩͽ�=�4���F �chI��.�>��<&靾]t弗n|>�~b���<��?�<�[K��:9=G�=�W��ې�u��v�R�����T���Q߾�� >�k�>e��=F�ؾ0Y��B�<�0�>׏R���<��>���>�4�9�摔��M>�/t���Y>�B>�ڝ<e��N>nd�2.>'����?%;l��>	��>5�Ľ7G׽'�J��F�T@%�8̓=��M>5�I��a�>�6�>a�E="�þR� >㢇�Q� =M>�ʠ>7х>�P>�\�>��=����=���o��X��=�B��o�A=�mܼ{h<<�����">��8>��j>��>7h�>K��=͟�;5�>e[������?���>���N�>Bv�>�X9�ǝS�Ŕݼ5�m�?H��&ϾTܨ�xy��������kk+�0\�>͙P>I����L>�%�=:HW>-5>>T@=�n>
}�<~X��Q�����������=��^=����� ��}��<Tݶ�������<6Y~>YF>V� >���>���>!X>VB��R<G^�>��#��C����ɜ>K�8�j����'�~sr>DL�=�����}=r�Y>���:i�=պ0����H��>"�>-/�5%?���`¸��*��#���]0�i1�{(��U��Jv<�5��0���|�<a��=>�@=����j�<�,%>�����G:~�9�Q⎽-��=�̽������T�<p�t�{���>��=Y[������<}�|�������kYT<1���Ε��į>�h�>�s>�ST>�%�>	�����Qb�?�,��Q�@�Ǒ_=�(�>ӽ�׼(vl�;0=ˢ����=<F��K�>��>�A>7�޾��>��н2�������v>r�x>�k�����)(�>���'��>cW�=�&N>T���ܙ�QV�c�5����d�<��>n&/��,>3��Bu3����=�o<?��?)��?6o?T:�=�1'���l[>�-^�j�=�
�>�=Ͼۆ�y��ߞվr�=r�kY��-�@>��Y���)�T�>,�?q�>��־�Xݾ=�>x �>� �>��@?@s�>o�|��0ż�px?&���!�> Ҽ,�۽�X��S{��ּV�C>�8��H��
O>���=þ��o9�sJ��uV�ΐ+�9<��y@7����>�&���W�;�u>��>�e�����k?h��>�	�>�}�>��˼ >y�>aS)>
�H�0L��$�O^�=� ɾ.Ʃ�ӛ���>a�W�*�E>`=u >:'�����3χ������M��w]�>�\�͆,>"�B��&�?^^?p�?~B?��?�G�r�f�&E��UT���Ȱ��煿m�׾c�d����R�}�־c�Ǿ�X��Q����-?f?U?���>��1?�<+?�b��Kr�=�X=��>y	����="�����V��н�n2=�8�>�<�=�d�%��>҅�>��3>8
�w�5>�e����0�����e=+��>l6��+�>3���̊�g����%�o�>v'-��Q��=$ ?u�?}��l�H��=�3k��`����c��f�>�7�=����@��K��i~����ݾھ�@=&M����tN�&�J>�_�C��>�z�>\�
?�߸=䣖��Ӱ�ߣ>n��?/������>B��>Se�t�۾�"ӽV�Z>��=?�V�=5*{����=��վE6��6��)@��G�'�Gs��_y=��Ͻ��>�Ɏ�<8���S'>q�>���~���K�8X�>ª�C|�>�]�>2/<?�l�>sY>�Rw>o*���bv=���=�1�<�9p�1�<������u�u��= ��>FQ?��_�>���=�)q���q���>&3�m|%>�!->嘷>ܟ�>�:����!�?�M?|��>�
?�֗>k���C>�>��|c�==r>N����T��鮎;���r#�C����;V#>>4X��2?@��=��a<��>��>AT>P\M��1??4����?�@Ͼ�[�>'�"���Z>����t龿����s����?�J�����>�Y&�+'>��>�y��դ��ARu?%A�>q�4>{��>���(��?�3=���)>kuj��5��&{��l�=��>5�y��냾�Lؾ�nA��"��]����!�e��ξ�������>�>��9�d�hg,?GǾB�>��讝�n�?���$�l(�%��=z$f�O,�>S)��r��N����>��+����ן���&>F��>�rx�.��<���>Ց�B۹>lS�>d�>t�>�i�=
w���C�b���9��f�w���=���S2�1���;�=v�<$_�=Zaƽ��>ر9���)����=~>}�1>��ͽVz����<3]?i�1>�!>3$?�=��F
���fϾ�ˏ��e[�xi
��w/�ـ>�7�(K>)2�UCI�cU5?s?ty�>S��>)��>������=��?���9�6"X>�o�>X9
?�da�3��>ю����V�\O;?��D?C(?]�	?B�=���`�S�;`a޽�ɔ�`C�<Q��=�u*>�����ݾ�w׽,d?9�>M>�>S�>\�Ǽ=\>h�>�Eg?f��>~�0�	����L�+�k�N�>,��=8��l;����l��?��B�@j��Td���X�����l4���������6֑�d*���">d6U��%�>a2��lγ�-^��@;|��>��<�H�?�B?�Z�>��S�`�Ӿ��?S戾5J(?�?�X��}`�q�9�\\1��@�=d�>��>�=~?Œ?$ >Rn�=��0���?g{����?m�M?��Ⱦ�ſ��W�������>Sf>�C8�������=y��xKx���<�^�>����$5���@ž���>R��=��>�|r>sM-=)�̡����	gK��%�=��i���Yd=�S뾌|�����զ>~]����>�=��l>0U㼭垿��>�=k6_���?
�:?0��>]�F>���t��>}&�>�K�>��%?�ٺ>l�7��+�>��=q��?���?o(a;K�>�Fj�	�?)�{��0?a��>K���F¾޵���Xݾ8�,>��=�(#����㖾�8��l���LR?rc?��d="�g�_Ǿ��>zf���S?�`?%g�>�e��V�Z߿:�� p/��[�<�H�>:F
����>��H�&=���>;4?y�>�%?7Xq���!�[���{�'�}>���E���Pž���z����y=(J~=Z���YM>Иɾs;2����l�=�B�>0�|��ɥ>���-���!��Z��>L�^�@P��+��<�-�>���>P���!����>�!3�޻|=�>�>�� ��WA?���>/U+>)4�j�?�i��]\?�\�#��$���e<�Ѐ�A'?XL�>�@|gC?��>#�>_ ���?B�=<?��J??kC��>W�F=�=��%>ֱ=��>F]�?mL�⭝>�[�>��6�@䡾�����^?T ?���>p����LGԾ�>T��W�=��8?�?P��>X��>@�1?6�?x8�>�>=y)?��?+�7?�U+?�R�>R��>:,>�w�=y�q4�>ե���F��?(��>B�w>X����,0?l�ɽy�G?��+��Gn>3:���
>�݂�~���"��l���)AҽPŬ>�]K=h<�e��X�>��p�І��h0��?�/����ा�>�Cl>��|<�{��:=��4>O�h?7%�?u_�>A/%>��3��8?yZ]�g�?���>�z�>�ѕ�<�ſv.�����a�3����>$o/�Ɏ>N�/��ޞ?S>� �>N�>�H�w8>�_�?�Z����>_�#>���=3#¾=0�:��>n�?�2�����t�>��̾G���Kx������L�����>�->yy>�B�t��=׆=U�عh�,��B��Y�>A"_��/Ⱦ��	��E��]����]>�\�1T��3�`�K�Ѽ�xݽЦ�=�~�>G��>#!�I1}?��m���@?�/'>/㖾�p�>zz<������:j���F;�ج?�ǭ:=@�>�پI>�J���Ӿ�;�,"���5>��}��m�?C,\>��=�5��D?�m����>OW��	�c��ҽG��� �v���=i�n�W���p?[ڋ>p�=�	��sU?r{�oY?�s��\��jk9��FH�L&
>��v��>��>eT�<wT����>�[>J��>A >�%F����>��V;Z�R�(c���.>�f�=}-D���/���.��G���d>�I�>�V�>�m>EG>�T���� �M$>�=�a�>��>Jٿ>�}�=#@W>MC�>��0>�×�2�g����C�d?�\?B^E�����ݳ��������P>Q���<hp�=c_�@J���>�B?�?�>��^����>?��>
n4?,Y>�?��!>39��;�>��m��`�=>���<OC��[�����ٮ>q�Yҿ>�"��4��Rt:?�n)?D!?��
?!,�>���=�/?7��>4F^�4VP>*�2��k�s�Q��%߽�ķ���n�&��L�%���Ǿ&ř�[�/>4@��i�?�I`>����-��|�Ѿ����Ŏ��Kr>��>�#�%5�k=���>��=
��;=���0C��/��b��>�H�<m�e<��#=׼�<#}���I�<�N��9.�����i��c����r𘾯���k%�O�O�墡=�=�M����y��=��ƽ�)"�� i?�Lľ�,>~�!? �)>��Y?ô'?h�D<�>�>�E8=Ӻ���?;�=�+��7>��>Qp��M��#�O��0Ƚo��=66�M8ؾ���<�� ��=Ӿ�~M���D��bԾ)�1=�@�ZT�>��8��Z�=��U�������'�<�H�=�L�\ �����z>�ܝ=����:��팾��>�Xm>��=S��<�[1?��Q?Z��> oֽm��=�}/=���=�]�fD>51�Z����i=8|�����G@��M���U���xG����/>�$=e�:�ǽ�|��_�> ���gƼ�=v�lIs>��>���>@
w>Ok�>9��>0�f>���ZQ���= J�>�f�>,n��w>xr=F͈>�܆��o�����#{��ȓ¾�!�wk��s����/e�}���L�=���=u%���DR��8�>��}>Ő>�z�a���a7;ݵ>�e�>�>>7��=�7>+�=&0�t.��3h=�w'>�T�D����_�>R��d��<Y�B>t'���.Z���>}���x��}���$Q��77)>
�ν#1�<�����>�]�>�^�=�~5>�V��!�T(��G��>fƾet����<�*���
��xr���VS�Q�B>��q�/yP�b���Cͽu��>���>�/�>�~�> D�=�-۽�ͽh�������T��|�N��d=u
�=���<�`�q$�QIp��\������`v=��rn���k��f�>���ӱt=IS=+ѽJ�>�>��>e!E>�ͽL}��?Z���R���>�+>>Eʽ�)>�> ]}>�"j�������:��e1�Ѫt�L�&��<=��	�q���=b�>uu��^��|��=E\�>p��=�ʾ���9j_=>���{~�U��>�|�>�����\��(�=�J�=�Ȑ>N��ے�R�F=�%�>�#.��^�7�A��4��7���7�\�u�"��9e�f�&=�%8>nm>►�]us=C9�>5W�>&��;�~(��^�<+x���|�(��>��>BYQ>�x�;P3�>�f0���]�$��;�m�>SI�����{	���>�=5���A������Z�=.N>:��>Jݽ9�<�rU>_��>��>��y=M" �go?���>*��>�M>�?Z�>{��>޽C>ON�>8	x�E7�=�F;���>����_����3>���=@A6<
�>���>���>�8�>YA?�� ?�ܼ�B>�@�< �>xTr�Vļ=#�a>�&2>��ǽr����ӽ΃c��Ce���T����Z����f��'���6=7)��3��dq=W�j>��>��i��n6=��>�T�>��,?J��>0�=����Ls����{
���=�� �,�R=�`��Le��rt����O�K���M�=��?1�?I<�>$	�I�=���UGd>��b��C��=�۔=�Ή�6�0���L�*�=�o��=���;V����J�>M�<�ho��׎�`W>�dd��m���ˉ�H5=���>�>�)'=��e>�F�>�~?Qd�>`�>%_-����Y��9pr>fvS�㭚=��=�.�>
�O��l�a�w�x�$�m9�<F����#=[�H>��<��k��8U�E�h=�k̽Y������oL<���>�D>�E�=Lc->���l� ��z���>!�N<75������@��+N>����Ž�<�s�����>x��>�?�>���>I�۾у�t︽�w�>|,��P�=��=�>2�=2��<F��=���<�9�>�}�>P�>�S�>��=Wy���"=�h">%_X>�V��.��N�<���=����}��pn=�?��>m�>b�>���>�o>o�>?:ѽ���.�<,q5�C�Q��{B=#�< ���{���ZƼ��r;��Ǿ��M}%�������,�F�"�'�o	�����={F����ؽ���Э�=�G>�+�S�@�۾��?�O?�C�>�"%�v�ؼő�=��>
5�=�$Q���j=�w�=+��=��m�]ᄾ/N�������t:?,?�L9>�s|��=�=�)l=�>�B>j��3p>\=��=�t��ZM���2���eR�>p]R<�����=mH>�� �A�׽i��M�t>��G����z��@��>S�y=��C>�>*�W>�3��4�ѽE<��"!>�I�[��H3J�4�V>�vS����8nh���>�">�[�=��=�9Ⱦ ]�.�w>{2�>�`�<�6�=���I�>��;>?>�4����>�?�g�>γ�>%��>�� ?w��>E�U>��ǽ�q>==��zw=�N=:C�g�==.T=�Y�>����������>~���|>���>���g�J���?���>��P>LeH��u�=��=�tc��F�>�+D�?����i=�!W=I���}־Ga[��z+>�.=��Y���=t!�=<	=)2F>٨d=��b;���>̳�>�{�>�m�>�����(���������;2���|۽s���J�S<%��
�+�	�"	�<i����q� �+�.���=�T�=2>ꁔ����~�L>RG>o��!�ϼ��e���>�PC>�4�=qi�=�R�=�|U�H�>p#�>��D>��A�su�=���=_Ο>��&�+UH;�ƶ=&��=sO뾮ۏ�V����J�� ?��/?���>��u=b}O>:>��F>�(>�_�<�̊>��?>ⷋ>��G���=2ʚ�������>+wg>!DJ�Ȯ���U<\zA>b�W>ˣʽC�=���=d��>��u�썾b�G��\h���U����>8�>!��>g�n>p?~�>�ӣ>���>+m?'-?﨏>���=��o>�r�>J_�>�3>(ڪ���>(�?rf�>I쳾57���ӽ���>8Ĕ�t'=uۭ=yA">$_����|��۾���m��H&c� DA��ē��, �A��=��0=(ֽc���% >W�`>FL_=Ӹ���^L��fH�sO/���!>��>�ֽ���G�>:F�>p�;cJj���ٺ�����z�\�%>�餾g�w�Ͻ�}�����ޅҾ�~���>M�:-�Ҽ���<]g�����=�X^��L��Vљ�7��>0+t>��|>F$>mD�>	J�>"��T��=<�>՞>�Sc�)�>�>`§>>�6�*$�K��tA˽��{� ܇��"��������'��N=C>�=�����v�L�=��#>\���2A̽2q�����Z�?�:%��!����\=��	_Ӿ��>��D>C�L>3ݾ��y=LĂ�il~>���觕�Z� ��t���ҽ�L��0�=��;>��
�.�ҾLrɽ9ݘ>�=s����\����W��!�>5Xv>��'>Rp<=�X���z�>��>5}�>D*���V���
���E=>;�?���><��=z4������Z��o��<�ꢽ���>��>�,%>ov���ō��iŽVV�=��%���@"�=G_��C��w���$v�d35��S}>�}X����ϝ���z-=kR�=��'=y��>�o;ן�3�ٽ���>��>�3�=~�>ç�>SE׾��ھ��=�H>)�q=KP�=���=/�>wĽQ��<��A|�>o�>���>>2�>���>(�$?a>�>�K�'u����=?�t>�\�=�U#�D�(>�F=��O>R,뾋�!��2�x��ղg�5�]�j��%Z���=;�5!@=S1�>oG_>�#5>}R�=go�> m�>";U>>�����=�=9��=������4��^;.>�����~<]߽,ȹ����=��������X��^Y>���>�}|>ˍy>�k�>½z>��>��E:��Q>V�q�&St�X���}�=l	о~K¾�t��m�	>�&�FRF��]�/IF>?d>�"|=����YW=��B;�i�����韟=Y�D=�;:>@&御ꁾސ���?�����ѥ�Sj˽�E�E�Q���Ͻe�=��=���=+M�����=^�p>���=qyc��^#����L�����Ǿ<��cH<���3�̾�g>oy�>Q��=����8��O�h=�D>�޾9��bq=�3Ƚ#?_��>�Ղ>7�>��>g�v�sL��o�f����>62��BtB��yO�9>;��=�f�<�C��O�Ʉƾ;�
�P˾�!m=uҦ�rP���缾��
>�26��������V�\>�)>��=.���<𿌿�����ZK���˽ǥ>�5>�m>6�%���3<?iQ=!�w��?���H�����>���>j�=SJ���\Ի���?_Ɲ>cN�=�����>p�?��>�὞`6��B��i�N5���G9>���>��,>��\?�k���Ҿr�?�ͮ��*��P�=�>?��Q?A�j?��<?sW?C���������2�Az"�[G�>�uj��ѽ>yk��⾑?&�=��B�e��6�e����Ji��x���L��xt�{a ���6�?f�=��K?�a���:]��ɾ��t�S�ڽ�P�b�x?��Z?ČS>���>F�>3�= WR>1�V=�[j;q�G��'>�{З<���=.sS� :K����>�����K��n��>2)�>�d5=�#�>�r�> ���u�є�a��÷>n ��3�>�,5?j�a?��?��^?)�R��v>:����-[=�~����o��'ݓ��~�f�+�+�Ѿ2�M�0U�>)���iY��9U����f�G?��I?�\���>&e�I���k�6'���v˼;����==�K4> M��qɾ]�O��{f:�����ڊ=�;���K��� > ^�>��>w������>�x[�^3-?�Y����)�	�?��#?^'C�Ee^>�z;f��;�;H�t<Dxξ4�9=��G�����&�< ?�a�=����p�þ6�r�%�q��6��W�V�',罙/$?X8�@%�>jA�[5��ԏ� ,쾛5�>M>�C�E����=B�c;Q���k�h��'�>#T�>̩=���_œ?5b�>��������U�S�q�׿`�
LH���e=����4��=zv���?u#���>��)���-��	h��r�>�x���NR��t>��W?Ͳ�s?N�>R��>�~>h�(?r=>sI�#u���?ߟo>�C�Z�=��L?�gվE������Oµ�-�v=�VϾa��>Gn�>8��>E�[�KZ�>�珽�93=@e��� ?n˄�,E��P�>�;�?�~?�>�6r?lxJ?u���dc6>g��ݑ?A3i>
х�T>�*K?]�ͽ�خ�g����r?;�;����>&��>j�1ɾ�O?ì?.L4>l����:��z?�$?��V��^Ͼ;k�=��F�%<{�L���E���@/�А	������>�z>�1/������R�^��񩀿|t�>�$�?5�=�+q>����x�]�#b��US5?麿��(u����	o-?,��>|񶼗纼� ʾ����EҾ*��^>w�=�/��t�}=i�=��>eo?��+?db����>O�?i
;?���;�2�>��<)���n�<�&w>x����	�>���@��=4�![�>Yß� &�<O��8�?�m=�3�=䕽��>CL�>�)?�?-?��r(>��h>�m�>*�����<�L�=C
?/AM���3������� >�j���>W��)}>��w�j���=����=�h�=�>��I���>���[�>�*�e>���>�R�=�O?I��>�2P�!2��2,���e�o�	> �w����;�$<�k#?
S#?�9!?��?x�t>*@��0�>��>�^���%����=�o�
9�>��4�z����>33�<4�>��??Ȯ�>	�1>vC1�P�	> �<1�K��K��K야�i4>P�H��;����>8� ?�~?�d>m�>�vl?�`>�WG��=��3 ?�i�Z���\����+iR��/p�Ѹ/���#�U��]f��Sb.��g��hn���JľnZ�H��?/�t>)�+>�ܽ|už9	�=��׾\�A���I?�>o�Q>O߾�?�𰘽 �Ǿd�����>�-�>�ݼ��*?+�*�?El?N�?�5�=6㎿�Q�#���^k�Krg��"�� ;}����>�g?%�>��`>h�!�Xk�>�0>\�������q�Y3b��!6�@��>-��=�����־�i�>}��EN�ڝ	�t+�>�B>���r��<�<�>��>ա��D��=�?	#>�2�R����=f�c�H:���ʩ�o��>��3�@�D��1���B�>�
�>�U	�5k'��|>n �>�M:���?���ھ�)-�1�?&����x��Ń���I>e �>oD?nv$?i�??욾�(6�e}��y�*�>�3/>r� �Bg�=��
=:Ȉ?B�>K� �`%��t/������N�=:�=�"�?Wc>�f>C���:���UM��������?��c>_�Q�E�W?�P��u4n?rz>ܮ�=z/0�Q�+>�?�f>ì<�TP�X���N�|�qO�>
/�bw��g�Ⱦ��[?�<$?�� ?J�?5l(�*���ы����>v���þ��������(>�\�= a�cz�E�?T�'>s!�=rX��vk����>趾�Ix?���=�f�>�=�8r?���=`� >����I?c*���C�,��>�"�?~n����X��C>Ù���ᔾF6�>"�>ga?����A�e��g\?3��>���d������g�J@�=L�w>��L�G��=�?��A?��>�L�>6k�@H.?7}8?ρ�>�!��P�߾����ؾ�Z��DӾw����n���6?E>��> f����?3��=��>�C�T���{��\�G�wS�>�j>�v�>�1�>��S?��?�6*?D�?�J'?�$p>�A@>��;)�u?��W?��d?J5?5(L��# ��eo>"�F�l����Q?�l�>uh~>�B�RԨ�1��>�Ĳ>U��/&	���g�>����ڊV��-'>�֗�m���Q�>���>4�Ͻ`X��G�!>A��=o�I����:��y��1ξ�����^0?�?����c>Ti����
=�t����"�?��>ҕT��[M?3b�	�m?�b�=BI�;��Ȼ�;���)�>N�>�����߾ϴl������]?[B�M�MVJ�7�1?.�?�^�><M�>H���Q3��w��D�M�r��>�C[>��?�\��Bs`?��>��=E�#�� .���� "Ѿԇ$���>��:<f�>���n��=k��<�>�M������2��$?���>��>Wd���})���n�Y@C>�l�?�M0<1@R���>	R=ԏ(���t�Ѣ�>��l�OT3��q����z��?\/?﮾�§�Jؠ�$�����E=U�=���>��>ڽĆr=��>M�T�f�?����0��	4?È�Q˾�e}�gDt�*�>Y�E�D[�>�Z�$֖��7?���>,>��Q;�q��4�W�L��4̾��e�7�ʾ�y�-�?7%Ӿ\��>� &��#F�Q�A?e�>W)>��=��A��X4�(|u�O@�=�����>��cJ
�1��>��>y>��!?&�2>Eg]�����_>~#޾����J��^O�=1`?r�>�f���>�mx>E.&�>l�>�ϼ=�����GS>�>�����	?:b>�>�/��K���1��o�?�˸>�:K?�!$��ae?�A�>��>ԛ��nо�:�]]=�eJ����A���>���=Jy���X?��	?.�9>W�ɽS�>���>�!�=�&��9<
kL?B�@?q�R>�������>E�L>���:�s�����d��>����F��=�>�X,?n�C?�5�?��P?,?s^c>��?Fx>�="xǽ�����`���{�>$+�>�*��<��<�A�>؀0�\�1�_	߾��?������j�q�!��kZ?iM����=
����gk���?�w��Niu���>�S��
�B��ݼ����C>�*��>�a��C|����>R!�>�?9�����=���=ٕ�>8O_���=??v�z�˧��X��``?ښ=B<��B���M?�O+�OS��"?��M?Z2X�J��� �3�>t(?S��>�݁?8�k>�B�>k0?�?:��=�L:�_@5=r~�>mД>�z>ۢ�>	Q'?�����\����=�jp�2ʾ\�=��n���=�"�h�q�.�3�Q?XSN���뾞���[Yu?_K>_L�΃�/�[̞<ҿ!=mt>4�?�?^˽Z�q�y?�=F^"�Ws.��Խ2�>l)c>E9=�-���4�=3n�;�=�Y�={8�<|"^>`P'>�	\=ĉ���k<�����=��0=z���`������� ���G�=�a���Ħh>`#��F��f%��.9>b�{�MI3�$���2>'SQ>ai�>��4>��>�X6<ې���������PN�=�q�<	:�0ɾ6ݰ=0z<��=#�0����� ���ν,ؠ�@�"��)S����R�5�;P�!@r���4���K�{�)�̽ơ�=89��@挾t�=�_�=d�>�V>��F>��q=@>_�=�f�/����,�=�	:���#��q	�� �=�4>�;s���>�>��=I�g<��Ľt���L
���fn��� ���<d^��hQ;a˽UN=�_q��,�>\>�9>[A�>�O�����Y���J�=-���3���9 �����g���`���,�p���/ϖ�8l�������n��7e>e@C>	8'>(&�>�-�=m�#�屮�X<�����1���D�i�>V���ͽ��=f����N=��h�|.�= =�H��R����E�=9J"=|H�<��н�n�=��/>��'>�(=6S->��I������1V�|ؘ�eI��uZ�=[:ƽ�6�w:F��� !$�~$��YϽ}=�6��;�tP�+ݽr��\���	S;��J���|=y�Q����'���[������.�G֨=�'>;���dP=W�x:1���;?����=[��=J��-Ƹ��x�=;[����<���R^��q��TԽ��(���%/�@$;����?���Mj�=�gνi倾E�<��= ����뽓
G=f�=0�i�����Q�j>Y&�=f`>���=t1�>�Uc�vi#�^���$Ì>G����ν B�~r�>.Y�xUν�ĽS�=��>��=2�>p@=�4���/�=���>Y�ὡ��+𸽸-�>�0h=L��=AN�=�a�>�O�<O>�=�F�=J�>�.ȽBJ<>t�<���=�Y����:�o�MLu>��*��RQ��=e #>�Խ�w>��z>�>���'[>��>��=8}��X:=NO,��J >.�~�<"�Q����F�������銾׎����m����<�9$<2w����p�z =��=.g�=�a����=��>�k6;;>�x=>��4>c�/����=9�~=UL��x��`B=ɬ���x�<��\���.��F�۾8^��aZ���q
>�e�=��q=�$)�k��=Q��=���=,�f�C��(��<%Ծ<�%���{��T�*��]�!�?>=n�=��>�,<�.W��DP�Mx?>��O����(>e.�<@�3�䪨��\>z}|��=qD,>��>ѫ-�uCԼ����t��=Խ�μ�R=��=ek��2x���r����<A>
0w=`��=S� >�Z��ks�A>�=�R�=S9���$������=� 7>٨�=&|=_��>�4>㍁:����D�s�->O�ּ���=�C�=J�>�ʯ=�%=��O=̎�>��>���>�r�>��>r5�:���Ѡx����==AB��Ua����=e�=���=�0=��=��>���>�q>3��>J��=������L^�=��=�����=ް4>�
��r*��J�"(=�[�>+[>HB0>U��>�T	�>�+��c=E�:!L>�����o佲����@�?��F=b�j�w/����~�OΔ��9}�>2������)��ҁӾV���)掽�2v�,=�������`ٽ�a��=�ʾE��=�� ������^������D��y��=���蠽�}�=!H�=-���A�"��T�=��=�1=I���ф���5��_��t$����5=:��=h�I���[݇=�`n=�Y�<�Ӽ�Ҽ��=Ev��,Ⱦ�욾Y]F�x���(�>�'�=P%z� �ʼ^i>�)�ʛ�<�8���l=�,����)`6�ߋD>1��=Is	> u�>�v>4Uj��˙��m�N�g=��ɽl�x�7Qp<�U�<ypF��Ƙ��Լ�].>f8=;R�=�9>'��<�\�oo�03��q���#�4�\�=N̽�h�|��<�=Ȍr>c��>]2�>�;>����5=$>��>����>�˼��=*�I��2�= B�=��=�v����ľL�f��&H�@�Ȼ�鼦�ݽf�ͼ�Ia���<M�"�-�W������fD=R��<	)�=R������㧻��=ǰ�=t�:=/�=�=ou0�(�U��<��=�O>��=�� =�v�=b;�>X�>��>�n�>�K���p��R����C���7��栽������S�9G��A߽�^T��q�<��Y�}q(�훾��;|�2>--�9�1R>2���ü1 ���>�"�:
g� �cf�=l�E= �=�1�FGC>sLI�;:=&5S=b�?�VJ۽�.�ک�u=�����Y$>Q�ܼ�A->ht�ݪ��g�d�У���1<ZA�=<P�=�{+>S�=��`>��;���=�\�=6	�;~��=�t>*MW�%����7��Hc+�
=��>�YS��yu=��=g��=��]�d��<ڤ=�G>^�)�k����Q���I�t�E���d>�PP>)��>�x@>!2�>i�{>v}�>�!?>���>ۡ�>"�>نm>� �>�̺>y_>3�b>�Rv���T=�Z"=�q��t�����=˯�=�	>h둾�,i=��=�w�=�ߚ��K{�X������XU��������\������E=6Q������vr=o�5>�?H=�%�����=�㡽h&���w����<:��<�n彙Q=���<���=��E��<{2�=q�>�{=1Ef�˅1��\;�&��^�=E��sЖ�Ƭ��˵�=][:�Z����ԫ=�{>��=峼�s#����>8Vp>�Vi>Pn>�!;�-<R�:�Ya��C>3]>I�0�6sH��T> J�=��=�1 �/<B���ٽ�<0Š�̟`�����07�P��?s�=�x>7��<3���Z��=rW/>M�=���ѓ�'>A�
>�ӽWH����=�0�= -��q'���=&#(=|�J>jF��P�P>�h/>:>=���0��<yͽ�9I>;M>*>��I�~=�>���<׼���t��Ƚ=<!<ؤ�V �<�>�� >#�=���f=�\�����=Ů>;��=��e�qa=��E�49>�>T��#=�f��|�=��j�l�!������(���g���p�S<�=h9=F(����[�<,b�=��]�螡=�%�=�i;Ò���AD�,{k��2��YV�;{`�<!Zu��F���I�<K�0�= W�<��=6��|�<f�=}M�>��A>Ypy>rH@>��L=��<lP��bE�=�R����+��x�=2�>TC/=ίI>s�r=Ʃ>�w�>ߞ�>���>Ȳ>�
>? >?�">�z|>ɲ="o�;��V��V�='��=�(>PɄ�ٳ}�a�����2����.������')��=���b���:�=�U�=F/�<# �<��>>� >�A�=���
��=h�=������=��̼6�R<0[<�*�=q	���G�=5��=��=�F��~Rn<���= ��>���>5�>�Z>U�>B�=vH[>�#P=-�>Ӡ!=Ǆ�jT�Z�B>(䴽8���Y�]>b���|�����Y��Pc��0½����U��=�x����(�;�D8=�j��Å=�/���EQ�N��D����ľG˽�$0��@�.�!����h��=�͊=an��݃�<Hl=>��
=i<d��.��=�����漈|���ѽ�殽\��M ���?�<�]�=���:��:>��,>��;.b���f=b��=%�=��>b��=�Xd>�>��>l�c=�
���&��Z�>�8�=�^�L0;]>�>���(k6������;��B����W��n����=����eG�����1��S�?��4x��b/�>hC;��M��ď��>?C1�2j�T�>�EӾg�ﾭQN�5������a�<*����Ǿ9�C��#�>�����?���>���>�2?*0?+�>
���OI+=�	u�a� ?w�=Ҭ�>؎�����#��VǾ�5�0υ�@�>�X�&k�>H}����⾿c[�S�o�����O%�>���>��?�M�>WH?�a�>���=*͜>h�x?{/�gߟ�$!?(�@?�D��+�>�$K>���� ��-�ݽ�Bq�̄=��3��)�N���~�õ���ok�w���ml����&�=�g�t
g?����V?�> ��Hk)?m[#�6�?�	����:>k�>=�6>(�0�¾�-��Q�*��n���W�M�x}d>�.I=�ʽt��\=�>/�����>�S�`M��S~��������UQ�>?E��y��>�w??��?��z?z�?�[y?1��?G����1Ӿ�p�=�;�?r��&���$����>$���4����\���/�?9��&�g>�m:��q`��?f^�>'�>���=ȵ �c��=�^�@I���w?*!��=�]��d�ԾM�����M������3?F)/����+1r?7庾�a�)r��t�i�?��bcc?�K��Qm�r/�=�4?��+>87`?��-�|) �p��$6��$>u:�>�hC?��=� ���a�M8>(��~FL���>>)D�����3�;�ؾ�J��̾����J5��
>��0�y��>��<�>��>�z�>O-�rt�>R�>�W&?R�	>��?!o��7��WI?8*?����G���w�@�:��ۼ����Հ~��!�?�*�S�뉾D�Bʾ&�DfJ>��H>�ɾ}��>x"Z?�("?9�$����K��Q��t����^?��?�`?��s?�c?�c�\՘>;�0����>
wx?�]a��>r��>H�	>U^�>��G=��>"i��P>�H?љ̾�i�>rq#��$?*u���K:��)�>�,�>���>*W�>im?~�?)�C?,tj��Y?`��>k���ͣ������@>p���,>��*���?M??���M��=x���>�����>�>��H<D0���7)?��=����FE��~(�?eY��P^�=<h���ľ�(�	�x��-�Tʅ��yZ�
�4�t U�݌ž9½���>�"���>K����^?Sߕ��v;?v�\�Ŵ�>yE<�&0? 8�?��G���=^XJ?"о����v�kQ��-����
��e����=W����W�쪳>x���C��>P"�=dc;���?���>Z�U?1q?�۞>`	/>K�?��U>�?#G��	��>$;���޾�汼�l>�U���S��V;��<�2�����Y�ӽA��=��&���	�d�>5Ax<�0S=󯯽�p>6A^?.������-	�_ܢ=��ǾQGE�6}v�2����U�C�3�v�>�Y���c�9�=A�`���52��!�f���Y������ >�e�I7n��i��9�z������ݓ��NF���9>��*�t���\���C�?J���E	<��>��0>�+���Ѐ>/b]?�E�>]�?*r�>���=T���x��/�������?��o���ƾ*�;>�������#h)?߄���	>���>O5{>h�X=�O4>!^<EȰ>�D#��U��8޾�`꾝O��*5=�a>y������=.�����>��?7�k��MT��?��>�Q>��\?���>X���Ѿ+$�>R��>��?�����?��E��:�=�6A���#�2��qNa�]r�>�겺k�d����������`>U��:�(�0�.�oA?��qr?�U�=Ҩ��h��?�x?o��>�٦=f�=qb�?)� >Qk�;���msҾ"V�`6��5�z�?L?f9?�q{?傇?�|��S�=?��/�z�>���>���=r^?�t��:o�^i�;|�3=n���,m��8�y�<������;��>���i=�6>��Z��
�Wɽ�`�<�͞���z=U�򽱊�=tp�~���
*=���d��B��Y�n��d�
����a�wx��Vղ>����Q>���>~��UD>���Ͽ>VҾ�I�ę���k!��X���Ӿ��8��>�*�/Y-��{|>vȁ�.T��[&>s�����=�|?c��>Qx=�����>\?��5�:b��������7}�򴀿C_���>�^+>��F?�7��;�??1R�>Qr4�%e:?�*�>�h�1��>'��=�̎?��0�D���"�A��=y�=3�?���o���
T�=w�^>;�?�����,��P>$��=#�?u+Q?�?��?���)���Ι<�����>�>�W�������L�>v�>�sξ�l����A�>�J�>���>�w �K�a>��,?��/�b<�>9�0�%�C?+ƚ�//V����>�q>72>a(�>9h??�?'�$�h0�>_�>ן>`� ���+?z��>{_?��T�H؝?����x0]=���Q��F��w������>���>��/?��?�?%��>[C�>���>�up?i`Q>�Q=�t��_w��(�V'-�1���D�پ��>>%3�?����K>�_1?�@?v,��r �>EН>�v�=�?���3�g#��R�����վ̖>�U�>�b{>���=�e>�CW?>�>���>ځ?�?�s:?#ّ��_?��>��>��ٻU�=���&?-������=ڋL�
Ƞ>�R�=_:�>�5��=�?��4�f>>ꢋ��J�>>t;�����ξ%dӾ_Ě�����9���W>m��=�X�����ݜ�>xO�>jѽf*W�����n�*����)�A�>�oI?�<=>$o>HC��i=s߹?ĐO>q`��'l.�WШ>�e>���v�a>.`~��������<�߇�N�4��o�呃���̾Ty������u��)V=��5>�!6?b"(?\��>��?�ҟ�����H�>0Ǿl���=�=�P?l2�l��>9��u�=&\�����;q�����7���-�m�fj�Z���>C>��T?yY��u�?�?Ke���x���,�>!��^���`v��߿�KD������-�=�4��/�>7�>��;�r��0��?�K����9?�o�����?�[����ZS?�#�KN����!?�b)�Y�q�%����9��e���6x�>��	��ݥ�ءn>�T�>�}�>EQ?/jþN}+?	�>�����*� �=�v;�0̦>�#$�$��>/����z���:��`>��6����`�=�˾I�>؟F�����Ŏ�>�#�=/�>�Ͼ`>z���^��$e<��^}�@1C�'���#?�2?�p���>X ?g�
?���>>V�>f5�>`�!�>3�6�a?�]?㝀>P >6����;�A���v^���>'ϻ�[����>	�"��;���M̾�B:������j�=�������=��<�)V?��D����=� �>�I�<oH�\��N�=&�߽�}W�@ ��w������+��P�>G�NI:> s=��?�`?�2;?�B?-�>��?�M?b?��?$?6?��\>�*����Z�j�	���Y���RѾ�������q_9��`�����53? �$?LQ�>�$?y?W7Y?�f?��K?��?\?��e=ޒ�Un�<���r�R>a��>�b0����;:���~\�=/�;>���V�>�6n���z?{	���V�]Ԫ�h��<:�.��N�>��L���z=}�?�O">�ZJ>�IV>��'���F��%�q>,�$���Ľ�G�>!��>_w*>�z&>��\?�О>�g>^C?����2�=*N��Z������tI�>��>�B*����=�Rv��B(?c�>A�	��R�>���>�Ϸ>�U�>�H�=�*ڽ'�?Z�=?3��?F"R?tqE?����B�>����t0�>4��>����1�=p�>��a=s�K��>&�Y�>���J�ὛQ���!/?a���z���O>o*?������ >��7 �?F�Z�cO�>�=7?����Ql>O@#��˿��L.�Kܿ���>�x4��b����!��?]���%)+>JǓ=�ŏ?)8�?�J�?�V?բD?�l\=���>�BC?H��4�?�Bj?!�׾_����h?�K�?&b>��>�Ҧ�)�>�����_���!>␉�W6���?G=ʿ�@	?B�>��j?³��-�V?��Ӿ�;=ٳ�?�xZ?�l>ע[>�s�>���>�lO=�L��Ⱦ�=�T?�DI??{������?a���k�����k��R
��j\�	�h�6���*ð���h��%��G�?���?�?�����>�U�5GH?��<��'��9P>+��?ֺ�6t����>>�D�>wjN���{>H�_>�����������u?3��>=���_���� � �N��?�A/?����_f�9z����=O9G?z�?��v?��?*�?�}�?u�������?}����4���J��w�>��c���澪�s>C󽌺f������GŻϠG>��>�wV�@��>t�>�>�>� ?��?83���!Ⱦݭ�>>�6?��ȾH�>�����/	0>;e@���=]��� �/"��F�\���?u6?f���D迊a��8m=ww?+}i?d�(?8��8��\!�>���y�?�C/?,���.`>B�t?p�?W��=�W�3oi�@��Hq��唚�l�ܼ�>?N�=�f��3jq��H���H>��e���|�lq���|���>�	��q}�?%����}�?����D�V>���>;1�>��`��j=�_&�������D&�>qh����r�&�t�t��>j
 �F�'>�ؾC�����ս�F�?8�=��>�܋�m�\?�|?4�?�u��؎7���A>�Fn?��t����?gTQ?t^?��=?^-�>>s�=��j=[&?H�Z>��3=�.>��Ϳ�% ?��ʿŲ��h��L@O�R�վ��?�?�o>��>,����ݧ=�Rc>]��)>>$�?�=��4�"?��>\Z?X*A>
��>Y,�=�M�՚�A{�>)�>�K�?����K�?�Ge/��L���,>��!�~�̿�(��;V? ��?iگ?;s���$��;d�>�3?=�q�?X%ݿ�W�?lR�>{�ﾔ1��1�E?g4��O�Z��u����z��U�3��[����p��"�|)��f#�>3ǁ?6�!?6�E�~�=ѳ�o
����?\5�>�c>xH��Լо�һ��<�/?�K
�O�(��ǿ�1̿ �?�v�>Gn���L���`>��3?.��?&�'�˷4��K�H�?�Z�>�YU=g�޾u=c�DC��l�>��;>�0?���}/��O*��Y?<9>ٵ�UO����A�>�A? �Z�E~>$ݾ������
��><�.?���>j}?TqJ>�U�?�a�$Ӣ�#L�>�̨>�y�>�?c�<f����)�F$�5S4�O1����dg>!V?���9���~?M����_���h@?�SG�/aG���t�\��^m较>G?@[���K���/���G=3b�����P�>/̬?Y�M�:�/�bB�fv�>]�&���^?]����r�e�9>x;�?��q�\�)7+�')P?�� ?��a�M?�����4�>�̽�_�?���>4�?��񽨂��E2>{ơ�ᚿ�E�=��y<7���3�=�������:*��0:?F+!�\~�>拶�e��=�R���=?4�>W$��х�ئ�?�G@�sz?jq�>Q���*>�)>�z?�S?�i��4꿊Y���G�>��*�}]?���=[2��'���c���C�a>��w�=�>�:?��¿Z�s�B«�� �?��� �ɿ���?��?��9��l�>H/�㝿�>��?7M>e,>H�=o\��E��F�j�2|H�3����B�#9�>?�>��>��Ŀ���?�R	����@�<?)�?�2?ʝO?&�>����[��ob<�s;�ie�qC>���>"�7�mE>�3>����D����W�V�B>iVC��������>6��=��D��lt7>K��<������x��n3B�8�=rFZ��)��?sH���?g��\Z>��>Db��\����?X�>	��8�ƿ�l=H�>�
��x~?��üsTi>�`��Os=�����>$˸?3�?Ź?���?SA��쬾���>�u)?��S>9�����u���^�B=��%w���R�:/��g�>'yC>�?'�i��8?���;F?䡋?GP�>�i�>���?[(?�q�޽?�[��K���x���R�c�A��U��'l?^M={1Z=	�?�k!�sP��h>P��?�a?>��?�U�?��e?�x��|�#\¾����CnF�D!����-?������>��M��i�<��|�̂y����=�ɂ>�>�=I�-�B(D���?�S?V���SS?D���Q�=��L>gB���ؿI�?����~>�и�潌?�!�>�p?\č>���>s���'�=K'T?sK;?���>�]>S�V?$c�>��a��l�>��K��3Q?s��>�u����>�.��<:��e�e/㼵p>�p����9������&��ڱ�k�������!�?��>�}�_�>�}s�>�������=A�ؾ%��>psg���>����mw�="s�*w{��<���x���?e{p?�T6�{hs?k>?7�5>��2>Y�?�O)?�B?Uc�>��.���y=�26>k��=�?���?���?߷�>!�]� .�>忾��??�rd����?C�=���������?���>�V�>E�=m��u����xA��ヾ��ؽ8��:�N����7��<q�8��L�=E[��s>3�j�Q �%<��ҿ�����?5;�?�y�? ?���2j7��s%?�Y�?�f�?:���05�m5�`���|��^4ҿM�T��t������=�zj��pF��/���R��T�>� �Mb�>\�b?�"?f��?��_?�UN=e�����>A0+>�*N?p����u:�dY�f�3�n��3��<���]�|��u���w�?<Ɯ�`>��r?[�=�����0�>�w?��=�mc�]?��.	�>Z����b���O�ŵ�d+m>=�>^M�>����t�?�l�?�G�=�����-?����:�?����m?�/�?#�\�Nڙ��6�?�n��W��S	���V��۽�զ\?�O%>�Ҁ�����%�B�B?�N�>I�#?=c�?pD���>��X�Oܒ?�]�ݰ��&Ȍ?X�|>���.��/�?
5�>@���y���)(�b_��n�o�~)?�D?�6�>Ra�@��QQ=���?����!��hF?H�C�4�˾����Ǿ�-��u�>2�?m_F?@��� <�	?t��>Ɖ�)�پ"]?t�'?��n>�^߾82�=J�5��>Z��>\�C�
�����>�u��->o�W?T�+>��Z�/�l>$QZ>��o	��?���=d���3?��>̫?��y��ֆ��9�>�ׯ? �>����>�5�=���>�k!����=���.�uc��e�7�� Q�7@�>BS羂UF?��y?P��>��?�#?��i>�w�>I��=�;�����uR=Y�?�a�'Π�7���*gA���>� J������8/�?:�x?�?/�?��?R��?]v�?��i?��Z?,=Z[E��¾�[?�x�>o�>�{�;O��>aó�q������h[/�d�?�>�R��&9��F»��:?w���ZK���x��4�� �>��{?����{4S��B��x?[��k��>��8>����fS�?̝�q�>P�E��i��
�?��>^��>�@��^�r?���>z!�=�Qn�C����ǽ�1�?�~
�n{��l2b��ɾ�x��fz?U��>ߤ��ꗿz;,?]O��J���p�����z?ɭ޾Ep�=T!?��f>��?�v�?����\U��Q�>Ul ?��y�����8��U
*?W?1���Jӿ�o�=8���ſK�ľ���?���z��}-��EV�>ߠ^����<��?.��?�I^��=�2?���=��5>��ɼ�~��o��gE��:�=!+�>c���=��ݾ���6��ݿ�a����5��u�?1�!?G��>S��>���>ؚD>�?��>u�>Z�?Z,�?}(q?��>��tQ=pz��_�#��⬽2�T>�$?�>���V��T,?���}���W�VU�>�{?��e>; #>�@$?R�>/�徉/���ka�ޗx�c(T��>>`9��xo?�;O>�4\��L ��)6>У>�G�>=���@�903��^��p1��_���f�<��bf>`��©t?���==w��ao���>�1�����>fr�WC���2}>��%>�0ξ��d�*� ��B�=�����ǽ��lj���{>�F�����Ĳн�X���g�鬴>E�>��'>��>9y|>��(�^C2?~�f�����H-���`B?��?E�a?�2_?۟H�iI�ԇ'�Gt�>jf�vY���ν��5>J������ɉ>�*?�ZW��=վ��k�Y���?T �=j�p��<�F��F���^�j���^2�y�"�u鉽CQm=�����=�3��YE���j>�^>��>Vǐ�Ǌ�������>��?�ҵ����>Tb=̂;��$?ˬ���&���1�Fd��E`=~�<E�˾�?1>��3��;����<��.>��~=�F��?Τ1=��>�?}X�V��
�u�J>�N�<
f���oi�|_}�?�>s��=�j��<�D�[>	�𾧞���W��;��>�h���9پ�Q���k��ml>|�=�l\���?�4?��b>�#��ɾ7���^��=F��u���r3E��0�Z�,��D���>FVq>�V߾�ԑ>��ܻ0��x�|m����p>m�X>�`轜��>�>���>��>x00?:*�=]�->�w=��o>o�*�WK־�=�=Y6?)�=sH�>�I���>Z�m=Fh�>k[q?-���+V>�`�> �?��?���L��!!7?������ʊr<g(?�ו>$_�ja��C�?r>>�z����k).?������=��?>'½2�>��	�zǄ�2>E&��l�?"�>���=Q���t�>0־� >ўξ���=���?h@j�*{*�v���ȡ��
�U����	�	�����4V���둾S'Y�k����>�%����!�=U�`��?�>J�?K����{�N�Y�u
����dچ>"�2��(�?�%O��=م�u~��1%��e+��쒿�R��j4?��'?Ge���Ǿ��>��X�A��<�Ω���y�v��?���?�H�����ݐ��r5� �D>69��������>Ê#��Q��H����>� o�XP����澡w�>�q<�y�=�௾�5>���>��g���!+>�U�E�<=	��	�D��랿�M����[?�\?���������Կ/ˬ��)��.�y��oξ�o>"��Z
J�	 ���X4>�+�o� ��P�0�>E��&н_���v=!���4U�#�{>�1?������>�l<ž~�>�@������|����>tZ?+?��?p��A �:"�=qM4?͵w��:�>����H����?�>� �stG��x=��y?ľ�?*fk?�6?iϽ�g!�&�C=�A�>p�">��s>��0��~���;ܽ�W��Ӿ�x�=k�?�k�>헩>�P�>��?A+�>�G=�V��E�?���>=�>	�ɻ���=]��=]�>���<%��uc�����/~/�ٮھ};�G����LS߾z�<�>->��Ѿ�&T?IP%�9�(�l��J�T�^��>�(������y?���>!ν��J����m=\z2� C��>����?�?�?.�?3|��E���|<��wQ�y�R?��>�t�����h�`>O��B:4>��0? cy����?���?��t>��~��O˾ա�4h����>vi�_���a�g>xi<���(^��,%�v�<�۾�	j�������g=�J���������=/�s��~佂�F>2m�>�2+��V�&~�_�>�����I0��&���:?�e>Yy�='d��6��y�{��p�>ڒ�>���>�]������\�>�bؿ�]�;��=�tS>�8�>��#?I��>]5$?)5?a�>�0�\�����;>m%�8�>v�d>aŤ��>�?�)~?�d�>jd`��"���h�V؇�h�>{�Η���#?Ӟ-?��g?𾣾�F �R�?HV���>G"�>=ۗ�gz�?h�W?D�>$*2������>���>.ϲ>q�?�,�>i�C>O 0?�x�eG�g�Ծy7u?H�p?v�k?A1�?A~0��
����u7 �����j>��>��1��zX?�վ<C:�K@���ـ�w?x>��>�o��p�>�Ă���`���3?�	��K���a�>t}>�3a>.d
��GU��r�>�!��J�`��~���M�>�b���8f?U��>��=��N�F-�>����1l�5��L)�<���?��{?�1\�Ԋ+��YO�V �0��?��?}V��@#�j��=l�j=���{e>٘W�.�~?p��?��'?�i��ka��Ӿ@�ݾ!�?������ <>:H�@���[1x>f�1?�@����?NՐ?%I�>��a�徔����2
��#�� ?�\]>���>�*?^�>�D?_>�?�/^>9)�?��%?5R�>//�>=EJ?�#k?��?��l?݂[���`?Y�>)hj<j�H�1x�=�^��Væ>:߾?�>�|��?��?��c������>�L�>�P2��!�����:������VG>X��;Ҡ��s�^��>��'>8u���E�RS�=if/=0�(�����'�6��>]��=�b!?�l?N6��q"��|�>���fz�>��?���@��?���>�J�>�,��z(�15=�U�>����X>/Е=�����>!��%׷�+/�utw?I8�=;�;�N�6��>�Lż��J�4�e�^E���s��g�>E���N�?3>�#>�&��A�'&<>Kü>&뾸_i�R$@�'����þQ&&>`�-��<���)��L����>��3���<�lԬ==g>�r>�q�<��+��ɀ�(M����c>�ա�[U>?�c'?���=���&��=��=��>�B���l��f��?��=?�C�>v��>x؀=��Խ��x��s��l�>��3?����N�?���=AĎ�VDy<z᰿)���O����?l�>�ʎ��*o��p���x���_��$O�G�u���,?�7�?1X�?im�49�b
˾��&��6$?O.�>�B��&��X�׼�v-�P)�=f��=�޾Ym�?ݚY?����󖲿.��M�C�=���>�����]Z�=dU��k��>��X?���>��?�m�;O�&>���>ޱ�=����?�W��e=�������>���>+�=�BU?����w�>������)�5�R>.*�>~�;?6o�>���>�1Z>\-?1p���龪�^�������<;R?-�~��?�Jz?�7?����@�=?߸>��P�[��(� �K</�K>
�C<)�'�7B?���>�v�>.�>'.?MD�>�	!>%Ji=kLB=L޲>w�\?W�W�D���>4�>��=g�>��.>�{��+?!�Y�����x!x��Sc?�?�\?�qA?>S?�f;?���>�CA�מ�>�|�?7�K�O=�(�=,�^��Mþ�O}��8>uEؾ�O.<h��e�,?ӷ�C�P�0M˾0�`��>�-s�=�)¾�I�?��\������J�6g���
���6��k$��p|>���=���=!=��(?.3>m#=��?��>�:D���|��̙>|�>��I>bW�6,�v�Tb�Ĺ�� �>t ?����<)�h�>v����]n�>O��ٽ��=�&?7f??b�>}?G=�v�=��(?���>��[��������>�g*��ȍ�Ί?���=��>.���M�>:;B�ߕ�q��z�>�eɾI�۽����XS�>��/��P;ڿ�s%?T�>��;���R�y>����6#Q�冻��E���ӽC�+?��ξX�����z�-�>�	���|$?��� ���m�?�f�?<L�?�?���?��?���RJ��A{?+�?j?�aɾ�!>|�?P��=
N�>����Ky>j���7�V?�x\��"�|d?���?��=��4>�,v��C?�B>Z�`?단?nH?;y�?@�?�����!	�@m�?RT�<�4M>�"�вU��an��1	>kNc�M��ũ��Wt���X������ʿ�sF���Ѿz��j�?�w7��G�?����O�?�Y�?�Ԛ>7z='*�?��R?~��>Uf�>��>�J�>ah�?gYȽ�|��Խ}x�>E�Ծ�nL��.��$�>�a}>)�hʌ���)?�*�r��� �X�~��>*�M��ɾꐾ"�\?$��>.�,?8�^��?����?�t�?�T?�i?���_v��#��������gĔ�B3����<�͇��ˮ�!&�=�=�̈́�|9��3	�Z����F?Nɔ>D��>�b����1������e�,?��?W����i��@�̾��I��ۿҫ��*F~� �����>z�>��>ŞX�t����>6�?j@�ܨ��p���S���m
��4�>�6?��к�i��5(>�H^���'�6�<?k=�H���P����?��?�*J?*����R?�-*?��p>��Ӿv�e�G�����w����?Ŵ��k]�/%=Z�>Τ��AJ�����2�?l�W?ݷ�<:��=Eˣ?��#?�ޓ?�5���T�?*��,��m��a=Q�~1(�Ĉ*>��J�=���T(�7Ć�=��F�پ�?�~���a0��W�?T3w?��R��WT��n�?d�?�?j!�=�?�u>��>
+�~u�?��?%����/?���?)E%�d�-?��T?��?��_�F���>���>q�Ҿ;�Z��#����	>�  �$�>}?����IȾ�`s�vVG? ���M1��l�>�9?�4?t,x>
F�>�Ӊ?�$?Q+?�eD>f�?�󙾀i�TZ?��2?�쉿�kE��-�<���>����|$׾�H�>�f�>`�����>q��?�z~>K施^d?��D?�b7=nJ)��ǁ�D���U��ó��c_p�kH��<�d��=����˿��>��L?~��zǹ��L?��>�	��8?f��"���a1㾽��>	K>АY���?
Y>�Q��@��-9?��.>'KԿlɢ�<Ӿ\���nJ���Ҿ�8�<�<l��H���C¾!�>��G��$@�QE�S�[���?6�μ�?�?�Wh�~�?��������>R��>>?q���'1�	�R?���?n>t�z�����>#�<>���K3���_�=qڏ����O1�I��=['��y?&T?N�T?��?{s������?08>YM����꾡�����>z�׾|g��@�C�d�=lF�6b��zu�S�>�K��:���9�>�vf>�ϩ>f͘>xg��|>��=��=�4=!F�>��ֿ�Y��d>�=Ez?��������{r�{	����L�+�?Z=��Q�(_�?���>��!?�Y0?����8�����>��c�a^�|���&F>�t"?�Zd���ؾy��=we�=��:?���>R��>W}��C]�맑�[/�>̷�[GQ��/}�-'z>Sں��\ݾ�(A��5����z\? ������={1��iV@G�k���������+�>��<>�~??���‾_־'$>8D�����\�<W�[��E�>dU�h����qY�G���>,�Y�W��ڵ>���?���Ý�*\�mU�<>;�����>r5��B�=W�?���>Ird�fʜ?��>^|?ҫ�����>��=�x6>z�>}Q����j��LZ��⇿s,@c�Ƽ��|���d��q��>��jE[?�oL>D�"?ߌ?��>+�ֽ�B&��� ��!��V ������\=�@7>�GL?�k����{�_"��e�>��'�hLD����XØ�ܝ��y�<2��>�LݼN�4?�f��}> (]?�C�>�Ȇ�+��1�>��>�+��^��i+)��D*?��l?v�>��>��N�~>o��?��*?ɧ��3�ʿ^`�=)�6>5��?�F?����u>?,nľ?3\輻�Z?�>�Gm?�@�?���N�N>�B �in�L�����a��p�����l�Ծ��%�=_����2vi�}�8?����;� >�C?
WT?A�p�A�d?�7-?#�~?)�S=�2�>����E%?NGU?�� >}�T�^8����>�+�?�?��Fi�L�ƾ��3?<X辩� ?)2�>�3D���>�:=���>�&>V���q���+�+�7�E�C���=����Ж��Ő?fÑ>���}ƾ!H���ν�k��p�=�����w�r��;��?����R�����6<X?c�����grŽIt�?����oI�=Jy >:��?q�b��?"z�?�h����SUO?!6?}/?�Q"����>JA�>)W�>�뽂���;��>Nc>�t��9�5?J�#?��>�[�>S��?_4�=�=� "�?�;>E������������>�<�˩����W?/:>b��>�Ϟ�oQ�>�V?^���B�3���S�z=�?=�T���`?����A���a������M�¼��>���>M�%?�k�>3�?ui�>��V?t��?t��=��G���?�,�?{�.?���>y3��M\�></�>Ieg�������?ٮ�>lN�>:����{��� ?��?�z����$>��~=�kK>�ھ`�>S$6�����k�=$�l?�P>R��R �=ڍ?��?����I��܋0=#�y>�'W���0>3?E��>�F������B@H�?pzx��^-?�w�>��Q>ݗ�?�	>�����f>�9�� "���/�.7��p*��%��ɓ��4C�!�<����Dp���j����+k?��?�`�?˵?��4?�X?�@<?�K���U�?�==?�D��E%���L[��IE�{���E3���ھ���>�:��[��6��lֳ>���=������=?r��>�ؠ?�������>���<�cԼ����U���p> ���ֆ�bbؿid�>l9��>�?	7����YE2?�R?�%п�3c>�nA?<�,?/��M�d>��ƾ�2�8�q�C?:@޾���qu�ANϿB��>���G�_�TB�>?�A���G�������Н��J���_�?M-�?��J���)�ss>9�>iA�>a ~�f̳����>�X�]x����>_5���6�����n?撗?r�q����t�o>���>�T��>�߾�lV?tڎ��X>�L���>&3\�:���ט?�}���:b?N�$�0u8?��O?*+�=ܴ��C�=zͱ>B����c1?2qݾ�Ð>@���Zӽ�
��K;�>6�B>3�����	?1V/���i�@�4>xv���(>�a��D��I��>N��>Y���u��{P?��>ȱ�������$?K?'6����W3�v�=�ق>�w*����(:��LE�B���;oq�-2ϼPM@?mf[>,�~>�_?�y?ҁW>ֹV���4?�@5?��>>���?e]�?m�3;�	�QP���[��C��:C���+�%�>� �>�.f?��?��@?�>6?y�?~�=?$>?~K?jJ�?��?���,2���c#?n^���>�>�?�c�>E����%�>��K�\z%��{�n 8���>⤿�Z8?s�%=��%�7��?� ��zl����l<�0\��7�?)uq��C���%�>2�(�����:+>ܲY?V	���z�<�?P.�?3XE?X=���
?�o�|g�?<4���6X?M_�>}|�|��<f�M�}�Ӿ����ր�#�����R?��i�z{ҾW�����U>1W�>�B^����3?G+��*9�?
 j?�v�?�K+=��Y��?�u��^e�>���>��>��n�����hT�>�&L>��>	����5����	?���у�&;��R���m���� �q�¾�
?/Q�����=C�?��?t�0XS���)�ܽ�>X���f1>��R���9<1;��߿���<�*!>J/۾�뇿�����T>��H�%&پ���`��?�?gp'?�Q�>`c�>X>?��>!v��h��>զ>1>��A�޼���O����b�KШ�L��
�}�8��*�y�,��T�>%Z=ǹ������!��4�>��?�k?c�A>�W�>ZN�> Z��?<Ј�Q�>�{P?%�Y�Oy��_�>��%?�u�=����?���|�T�L5����C1%�f��eX,�ѵJ�R0�9���T>;Q����n����>�F>��ھV������>P�>W��>t��=��4>��>��>���<d�OY��,�J>!$W�P�oK>��>�-w>cU>��̼�N��h/�,w�˸��M�q>�>���+�N"�>Q��>=����^����?��>?�?��>s_�����]�̾�MA�6�9�&X�wlU�a�<J�v� Ͼp�j:��O�]![�Y�|��e���u=���>B{�>��%���=tE=>_���M�=��7�k>���ݣ��e��O׶>�ξmQ��Ro>�@?�rm�a��>�\̾���=����z��ѡ̾�	�>x�t�1t@��ݙ>��>�i0��n!�$G����V>UN��F�>�񎾿��=�F�<�0=�]�>�����v?�H�<�?�=����-c�>��>����N��^��Y���]��<�R|>*����E>w:�ӡ�>ʕ#>��>	FE��?9��>k��Wf?LM�>To�>i�>�N0>9!\?]B�=��=D�/>%V?��%?��dɾ��c�=4���=���*���3>e=|�W��>7?���,M?BG>	�>m��>���>�l�=\�T�p�K?��׽R��Ѭ]?}�M>i��>�e���?��W=�ۖ��g >_�u>Zl���򗨾�>J�=��r�׾0����>:���s?�k�J�=�����>	_T=)h`�۔
>C��>� �*�=�X����? =�>��I3�>ud>�]�4m�>�?���>u�
����� �\а>��׼L�"�C�>�)�>���G�?3d�>��>_#��"��=��?ϑ?��;=Ԣ>/>?��> {>�D��]U>��!?�te������,�u} ��3
�j��ٜp>�C;�㾑��;��X>���=ڹ8�\�Y�:­=�\?��+?�t>�5?4� >�3-?k�>�߀�x]S�t4?�O���?��B������r��_��ھ�����M>n.�>z��=��"�)�lD�>�W}?����9��1Z?�Z�>���Ҍ=���=����9�_�[湽�-�eH>g�������=�3>�?��I���u<�x���N>yb�6�=�>1e<KEE>��)>��!?�;j��@��CH�<G=�=�QF�X�;�iLԾZ�1=Y ����L��4�C�>���=!�V��z>_�X>�8�>"��YZ=��>R^�<c�;�Q	�#<�=2?�,����=pʨ>�"�����V���ƾ��>Ə̾Kf���>�Nz>���]�ؾ�����>ng?���>Ce�>��Q�dcþ� u� ��S`y> Ծ�u��8��>Ƥ>9��+>w��3�$?"0?> ?	�?��Z=��e��+�=$�=�*?�����>�?�>�E�>����ԾrH�\O�>(f�>��>�Vl>I �>}ȧ>"�3>�s���f��-ٽ���=�\t��a�>'$<��̖{��d@��o����G�~ξbw�5J���_ ��\��C�>��ƾ��L�n�پ���>4ů� ��>�#�S-�-PM?о��~�+��%�>t^?O�>UF�>%�1��$<?)��?Cv��P�rXL?6��>���>A�����:�ᰢ����.��>��>�>e?������>�3W?��d����,�>]d>�q�>�$�����!QO)�'[;>��o��v���I���>��>z��Sݱ���!>k�B����[����s>�L�>�ݼ��T�ry>Oލ��mq��+����?4�6>\� �x�&�4��>��սƝܾ����?�>�j;q|�=s��$��j��r	��*��jG�UM3>~�=	h���B0��;�J�>(�>~I�>РR>p-�>-.�>���>�b>Я0>��+��j	?Ge�>kȾ������?	�H>p��=��
�H��
�:�
�� �d,?Π��~I*?�'u>i�=?�B\>7	?A�1=8��>��g?h�f��_�����>ܿ?o�7?�����Pc����Vy����<��Z�}���s^>14�>�)Ҿ��> ��=F��>�2+?w�>��>�ܾ�����D'���=h����F��.���s>���|�0>��&�H9�>�S?F�ܾ�%�#�8����>�60�cL�>C���\��q��� �k�3�MR���o@��S>�u�<�ҾT����>�<��u�>��>(�>�����b����?��d?-�Ͼ�j�>�>�fk>F�����f�O�.>Ж�=~\�>97�>�[�=�h>~?�����>DG?�ʽ�U��e�7?sć='���#��qiϾ����N��aJ>Fm�>��>W�)=��@?�PQ?\���u�����A?��>�p7?�R����Վ�ڛH�Emᾞ; ?��_>2�?<k�>��%?9	�>��h?��?:SE?�	�>4pG?#��>���>��m?bk�>�>�>�6����;���>��=q�H� �F�Zd�>ZC�?S����;=��>M!�>~�
��+�0$>���=�1
����Ԗ�����Bq��w�:����Ա=pU����u>G��>߼��������� ���� �^�-�\N�>�t����>����.?e��8��>4�u�aS?W�/?O����Ჾq>���>��>�S�<2R���0�C'�Kف>f� ��ZY���q�N�t>�I�(��8~�<��>�I�>O|�>�<�>PI�>�a�=�f?���D?h�c?��<�bV��H�>�Z?Rd>5u�h؝<K���:K<��̾����+���7<,ʬ�%��=���;�9:>����l�<��'?���Iռ9��#�}>�����w��Cb��7���>��龯�1����< s�>� @=�<�{�>AՓ>;�&?����Z��K�>���>�s?	�¾��;>5����1��?��j0B���tz�>_ج�a�D��#>���=�b��~�8�����p��V�,�>+.���!������>��f?d<G�5�n		?���>�"�lK��剾AZ#�ґ�`�	>��:>�3�~�D��׽�2>�#K?1�ݾ������>�^>˚��_׾��u�{���m�>���>�5?ND�>��>ꥮ�BZ�>�g? �.� MO>4�>eג=*��>��>��*>�&.�!ߙ�F2U>���=�|>`Ȓ��?�zK>Izp�H��<�t>=>f$�>���>�W�=^:">o��>e:>5C|>�M཰�=?�~?JOþ�{����V?�ܕ>__N=;��Fq.��Ѥ�>-���9�I���N{s����Yw�=I���X�=��X>+��>�����L>�'?�3)?}M�'�4�<l.?	�b��BN�|ϩ�p����i�x>n�:�	��^�>S�x>�����0�ef���p�>�4?��?��>Œ?8=�>�<�>øq�F�>����j⽷׀>�ft>/�ֻ�@	�����f�>��"��	�'C���N�>=Rw>=:a�L���x
?j+;�-�r����?b�B���K�w!��@����~����!�4���g���<��ƾ�V-=���=��>"�ܾs�>	�2?���Aw���?��e}>C������h.��H>烅=ٜ��K��=�?Z?�"�=����	e?�9C?�VP?�������Ø?H?FA8?�[�>?͡�>	�*?���=�M���?
�>ޞ2��^;p$����?�%׽�YR�H���C�k��8h�l�ԭ=m�+�D�<\#��U>Xb���NN�.ɾ6>JX>��	�,�����P����m?�?�?�
�R��>��)>^�ܿw��2a?b]̾(.�>
��<8�ٽ�����Z=�:�?��>��>E�D?�y�>��K=Ќ�?x﻾>G쾝��<�Ua���2�����-b�G��ر[�n��>��ž/K"<���=��"�"��O�>\b˾�n�;��?֒�D�n=#é>v��>���=���?�
�=��w?����0��NE�>� m>�uT=���p_>_T?�I�>�����)?h�C>R_�g����������z-y�r���Z���im�y�>[EP�_��?��۾t����D��zm@+Z�?zx�?���?%n�>�D���R?6ڤ>r�о<�@�'�F���]�&_�� nZ���e�!<�tU���X=n��M��2!c�:��u��}������;��m����>�֓?�cF?��>�D�?�D[?K�?VV�?hCv�:���?%�=����{r?¬۾�h?�`,?���>���֟ ?��e9Ҿ���F�/?�C��{�T������9�*����k��Z��h�>Ǜ�2s>�@HҾ3��>���)�����j��ҙ��a���C���<>e�?���>̣���o\>&瓿�$?�3�>	��ĊC?�����`�X'��b�=Ǻ{��������2U��N���Dh�>�ľ+lѾkUR>?�#�?n�=a��>YE�>���>@�q���I���X���h����U�[۵>�;��x[7;!X��'˞��vT>�	=?���=�ʹ?	-�?I`���0�-@�?,T ?�O�?Nc?�l�?���>��>�%�=�?TM��s ��թ̽M����O��Oj>`0>��\�w�=��+?�+>���֬�>�
�=���>��e>l���>nx=��?���?��f?=,?�R>�-?Ϟ�?���>��O=�ӎ�/�/�*��>f�>,?p�O?_F�>��>��?NV��ǐ�M�>�|Z��PM~?Q��>�`�>1�?Ec�?�瘾 ,����`�&?T�>V�?8\L���?o�ϼ���>���>]�>��w��ܼ>ug�.@�E#�J_�?ĕ�����>z�����J�*�8�?�l>=����뾮�'�]�>�4�?��ܾ��=�n��-�?1�0���>���q�>ɿļ��^1�=%�>�m��]�U���o#\��}X>�#��R;r���?��f��+�>/����y�?R?��?���=�a��ýB?��>9��>=7i�
Lk>��%��D��7��~�>�����>����5X��/��"���:�?��.;��#�2��=�Yf?0\�0�?)��ٻ{?|9�?�n�>�ӱ���$�K鎾ɨ�ǔ��]';�����>D�	�OC����l�V�ھ*�1��MK�������
>��9?G>��Ŀ�>[U�=�a>?u�M��c�=U?� �>.�'>�-�=��?Q==Ҁ�>��E��-��C�D��6\��m3>�9ľ���pT�1��'<��!3>A�5�:���f8^�B��O�c=jA��T6�.�ʾ�˫>��6�A�?�P��w���~����3��J�?�:��p)|>����i6�����C�R�>r�P���%?;��?�B,�^vx>��?����;)?��E������?�TM�gd��A��M?w<a?t]�>��+=�� ?lN��ͣ�(�1? ��>3��b�f�L;k��l���1���+�9�ݾ1H�s�>&��&���hZ&?���U�>5�?C�|>1u���h9��$ҿ�q!��Qp����>�8G�K��n�G�0�����pd�,9=�CX��m���־'�>f(��u	����Nm�=��ʬ�=���>Y"�>�t=>����h ?@�&?)�=�߯�5	~=��?�>�?P��?��!=��>�d���S���༆�ܿw��������>��xЏ?i�6?�S?��]?��>��;�?�B��}r����)?���>r��>���>܈Ծ�.�]N���J?�7-�n*\��|>eR�Mm������n��4���z������^s�>�Q;���>]��̓ �x�_��u��ͯ��ℾZ�!�B�f��J�e�h�(�ÿ���0�$�?NZ̾)�Ѿ�Vӽ/G.?�½㡛�Y���,I?�N��Hl�>	���q(���lϾ�]I?2o8=�^Խ�>
��h�f��!��Ș�<��>Vt�?~9;z�?�F?�[f?Z[�?�P�=
��:�˿�A���K�<��R�L?xO��*�>�@#�쌽?F��=3��==F.?:��>D�?���?�V?H_���XZ���>������=>DF�d���5�J�c�?�m?����>*�E>wn羸Y@��>��4>�<d?���?h�0������> �1>�� ���HJ�=�9�3���@��?�����+?��?��-��WC>� $�C>�d?�+�?�4?��8?==?���?�/�au���
��i?q|;���>��ǿ!G�?�=���?T�?�E?#�B?���`v�>q�=�O�>7��n�?�
,?>�>�
�;��ھB(^�&'��˃��ʾ�!a?1�?8�?��@�}?��?�?>�~���Iɿ�����]�������}��>�?>�ǜ��a���g=?x��>ma;?�I��	��>(J�?�Na�`����>���>?��G
 ��lw=Hlo?~��3H�>�i�=U?��>թ?y�*?��>k�?<�?�BP?>+3?H]*>��^����=����<?�\81��{=|�>����̂ľP��?�
+�hsu<�F��,$>ӽ���'�<�W+��KR��8T�%�о5�۾s G?��>P��01?	��>�n?�� >�0������i�ʙ�����=�]�>���>	���\�־��x�=>+YP?�s>��>�6�?�E����?��7��=�P?"��>��p>���=k������#Ӿ��_���:*d��N���#�>7we>��@��\?hi�?�
@�|��(xʿ���?9陿���?�-�?�o>����p[?��0?�Q=���v�*�ғ=GE�;�ʾ<���A�6AN�[�]�R�>B��>�,�=A&����*?�����?�~�>`U!>;�>S-�?��!>����vI>�(���E��U=�Z#8?�-!�R����J�Y��?[<A=H-�?��vi�?��ݱ�>��J�B�c��=>��?� I�#�>	ʖ>�u��׋�=@
?Wt"�
'�>p���|�X%i��OŽOa��|�?_��>Rw?GC�>%u��j$�<�&�>~5?6�g��)!�@Z>ǒ�>閅?����BE�ڟ9�h�>I�?��/��m1?U�+��R��{D�>7�?����ľZ_>2�y?�פ�궾y�=9��?i->~�~�%�þa�;8醽�l�?���>"��=�@�>�#J>(�չ���>v�k�����/����>�1�>��<��Բ>�9?�j�>3/�>���_��vZ?���>��?YNk>ެ�?.�a���?s!�����������	��~�>�z�>���>#޽�z4�RS����p?&�H�ʱ���H�r�.>��¿�N??��վ0�g��%�>#�(�u�?Y%���>$��?0�?�����?)*۾a\`?Dm�>d�w>Q�>��B>����I�>��ݿ�|�>��8>��/����,H�v�?7�H?�?]bW?jr?���>�颾N徺E�=��?+~;�Bb��VCe�'�<J�a�F����>?�aO��=6����p��?EZ��$��Ƶl���?v%=��o=*��>�8?�m��@>�>��;�39�?����B_ ��r�����$>p�r?�K�����?2��=�(>��L?|����h�>���=lh?.AK>*���)&?�+���]��=�\콴�D��eM�����y���,�!8��/��nJ?�)ӿ��@#	�1��>�z��i�=J�=�ߗ�dm@?;?j�5?،�>}��>����s���x�>pku��Ç�D5�=A��=l᷾��+?1�N?Z��[:ξM{@>l"O?@=�>���u��Ó��d?VCz?��ſ�'?�2�=�5=@s�*�V)�?��?L�q=�6l=8���=H<X=/�z��е�����,h��_� �����#b����=����џ�:�17=�/>��'>���=�`�=���=+=��'>�F�<�� >��=DO>ڧ��I�!��5����XAk���!	%����<��+>�ۂ�G�=��G�Vdv>�yt�< �;N������>Ԓ�=�T7>��e>}b�>f�=[��=?=���l��(�����=�<[�����=Uon=7��=��S�3k�;�OP�q�ڽ�6^��}��]~`�ο[�7G\�=ˊ�i^���R!=�h�=�<LS>tѽ^]��_?8>����(�ս�I>`[�=�=��P=�(�=U+���EH�S&o����=�]+�71��2 =��>���<�aP=XuS>[TT��h	�|���ڌ=���ֻ�!>w��=�S���#����)=,Ҧ>��>�X�>4С>?�q����	}���{���
���作����ͽ�uc�]洽q�w����L���N��´��>���b��=�.p>	��>���>�(�<�t������+�ļVW�=�M�%S*�g������fr8�,i	==ke<���:������<e�3>Fd3>C�����<�)�=��_1�I��<��=���=Q��<�1>!��=��9����,ݽ�g��]u�=Bi�<d�=��Ƚ?�;���<!b:;cG���tӼ�X;��>9����3]�e4W�顜����b:�Ŕ��_=�:�G�+<m>}�$<��㽪�z=��X�]��<]�%���n�8B�=ԶԹ�5{�.��=w���
��v"�jJ%=�o��~c~=>�-�S�)�v�����m��k���LO��_e�����xg�\���/>�6�<8":�Q�</K>	��=������Y=��=Z�M�g�6>��>c8>ϭS=�K(>��=ʹ�������>��4D=�Q��<�L>�\��P�j��5�<���<
3Ӽ��:=y
�>����7q<R�F�>�M=�}�=�*��>Ś��J=���=".�>zi>��C=H�=Zv�>
� ��rI�1�L�>E���@�/=�	����3>�BԼ�m���=��㮙>k�s�O�Z>h��>Ֆ�=b���Te>jƲ=�*%>Q@�ɉ6=E�>�!W>5���&Q�,��G�[���?���$����w��Y���M��g��m�=���Gc=8C>�\b��kc�8��=r��=��<F8t>���=� �<_�p�Y�Ub<�}���a��^#>(g�uH2��e�#2l�{���j�M��0�D����-��=��<R-k����=��G>�[a<�9>��\�;ғ�<0�J�{�r��"�R�	�[����<>-;��=l#�>�&�K�溭<R�>h&=�a8������t>��=�1�=���=ɰ�>�6>�O�=��>��>&�N<)�I�~����xC=֪�n�������跼BH/�Y�a��O1�v`Q��w>R\���M�=���=xd�����!=6&`=*ҽs� �����]r>�t�=�V�=��>��>J��=�}������o�P�=k�<=@������<%�c�����;��=�ͨ>�R>?�>�m�>3�@=����*6��n=q��f�H�#V��3>o�8<�*��W=ђ>^��>6O�>�W�>�y�>�}0>�����;���}�=x��:G�*���=���=�^=�mK�*:5��.�=ң>��>⁙>��>��F=��	>���>��<���=J��<.*X;�,۽�	�=�5=�}3=DAݽ��׻���XrS�O�N�/���K�p��)�Wb��3��k>�I���}�X�">UG��)nI���r���L=~�=D���l=��g�R�
�0>����,=�6T>�<��3���=��N�Z�>u�=��=�ו�f����-�,׃�����«�=�9�<�=���50�9��Ӽ�'�<�o���H�=1[#=h��:����r���h���p��QG�>�
�=SL�<>E���4">5�� �@�η:�;�~>��iwd�5��0Շ>��=���;��>�2O>z�V=�ֽn��r�=���g۽��M�>C�5��~�+݊�E)�>�i�=�Z={>>gh⼬�<���^=�D�=̩<���=K͈����>dT����<�=���>�mY>�>�~�>� �>ؕ���=3z��_es����=�@�Q�ؼ�d�������=��뼻9�;���\�������ʾN1 �9�ɽ��}�˽�5���"~=�-��f)Լ�o��>�����/�`-�=�y���_>����TҼ�ъ���D�!,Y=��_�O�(�N>��*=��=��v<��潗���%����u>�#h>"�>QƩ>�ƾ����?��>N��Z�L��e�����¾��@=z�Hw���Y�G�m�^�:�N������#G=��Ҭ<�ϙ>=#�3F�9���m�u>��f=�٭��Y����=�Џ�˴2�`*�='vH>����y*-=� �<[��<�S`��wY=t��=�أ=��4�X?>���=.��=�-��F�7��y"�e^!���=�9>�7=�#=�3v>�<ڇ=.4�=�ݼ��=���b�=5@���*��� �M��j��<lz�=�:���W��$���Q >\b�,P���˶=���;��=�逾ƒ��v}��j��菫�Ĭ�=F>F�:>�{>f9�>�u�><ނ>�-�=��>S�.>�Tp>[�D>T�[>��>�J�>���>jۖ���= @">�F��~�G�O�>
��=�v6>M�����=�>:a,>򩛾��_��z��ܭ��24��1��*��,�a�s�Y�==(�=�y����W�=N]�=�[7<�s����;ɖ�
4��w�G�<��= � �9}���Z>ې��&�=���=�$������=	��o0��E��+p< �{a�߸?��Ͻ�k��Z��=]9��^�;��>=قe�iaн��ֽ�:>�o>��v>�\6>�M|=x�>���<
恾���<C�c=~>䀡�ʫ���='9>��/�ςͺh7~;X�2�Km��=����;9�h�l=�G�;=��>"O<�yC�c'^��)C>�5�;.rƽ�u���<��=Uv�Ĝ������Z=�A>SDi�u'P�F�	>p �=w婾i&=4��=2D�<7M��4ؔ�y�=����W>�po=���=��G>�@=�9ʽ~�n%>/a7����;Ma�=��6u�;�L��5�=f�=��b�,g �m�+>���:Vτ���>�:*;ڈ=ַ����a��Ə=I�����z��{ �A��W�\��
����<�p�<:�����|�2�_=��[�0�<�a����=bS�=�A�v茶�"���ҍ�p������A�߽@��=���=���EMe�Y�=r��=�=Nd3;�ܼ���=r�>5y>%`@>�c�>z>咔���y; ��=q̉=ˣ�=V >�Z�>��=A�V��?�=N�e>'�p>�n�>��_>P�v>��2>J>�&Q>"�߽�=Y�>��P>�U=�箉>(��=ro�=ax������t&T���A��<I�S�k��w佱�������N���=3�>�W�=8\��A�}>B�
>��L=R�ܽ!7!�q�<h���}
>�l.���<_�c=qR�Gn��*��=���<|�=���=��>r~�>ƫ�>���>Ӥ�>^�>�9->UF9>k��=D�Q>(TL��t�ۗ��Y	�>��Ƚ�~�G=nB&>7�˽D���\�=���4� ��b��ҍ�'@潩/"�Y�t������ȍ=+lw�Ar�<+(��9e�FG����X+����-��Z)��hF��н�m��=(�=�J ������޼	*�=�>���=��9~��9�����-������,O��nĽb��NiļƉϼ�v��k���?<>�h�=��#��I����	�l�;�;H�I�>�\>b L>�~>I�>":#���=y$�?؜>�ŽD�;O&=`�>��;��r=��=B���3c#�����`���^��x�9�����h���+>]m��Z��p~�G��=Iμ'\d�!F��ޟ�>3�?�T?��=鋴>�H�=f�'����?�':?�Vu?�����I> ��<���E�[=��s?u�D?��?�E�>g����c�=N��:ս��>?��b���l���/<�����~���`@�N���L���W�g{.>�A���'3?E�v��ڤ:iС�'�a>���>���?Ĵ(��k�?���?�e/?t8?�E�?o�?C��l��Ͼ��9=8/7>�W��hK��p��Ś>���?�D;%�7>MP ��{>5�վ{ې��@���#轧�����.��?%1`?]��>GẾ:>�N�?]E�<Ɂ�8��>�b??��=O�?���>�QY?>��?� ��ߖ��w��� <�ǐ>��O��;��7q���:?�(>�/���� �H���Ͽl��_F~��Y����>p���ھQ�`?2?��q���A(�o0K?�Sg?Ae?�?AU�>o�E�g;#?S
<�TQ>���＾=��7?�Y�>S��)���>�ā����>?9'?̲$�z�z�O?�O����,�"����F��7����>{��>���>�&6?������3��6S�r�9?�L�?`q>�<���B�������׌�bN�?����7��=�K]�J5?�:��ad���Q������-�0/�=A���*�I z?�qj=�w�H���o?%�?�Ǩ��J1��@��ܪ߼%���ɬ>~� ����>�{������&?�Q�>~�e>�о�o����>:wO>�ڗ�L6z��R����=f?l&3>@�K?�?�>_4�:>:�����+�>�I���>
�n����M�E']�'�n������Z�/Z��8|��l�>~�U?
IL>��a��sQ��>��h��U?h����7���=K�?�yL�uŽ\8����>�n?=�<?��Y?AK?:2?�c��>��<��7��?	R��Hb/��&X>�p�>\E?��Qݿ�,>Ɣ����? �M+>Q~����f>�� >7�>�zҿk4o?q0�?s��>7䎿-�?X>��Z>z?:&��M�@̃?rI3�a��>�<(��!>	&�=�3d>ґ�>Y^�>���>��=�@�*?���?��#?���B�>�?�f9?��AV)?��1?l����	�T}w���h?��<c�����L>�?s���Է#�Z?x���^=��>7�g?n��?nI?��>?rcZ?��3?�A?��J?��>�nR?�Z6��x�>����-?9%�>�bb>No����a{����������?a�����>g�=�Ψ>kQ7�������&?A�A��NZ?2Ͻf�G��$�����@پ�`?��(��^�����Pi���H?y��=�K���-N=Rq�Zp��Yb�>�_M?����?���?���=VR����?�?|6U?�`�?G�#=�4�������=�*�>����ء��-*��"e=���1S��E��%0����@��>p��?�3�?�5.��ـ?�0�>䆽�	�=�O�?�4,��A#�"��>Pg�>�=]��"ž��>��ؾe�>��?��ռW��?�w>?�۾R9�=ڴ��������>�ߒ?yH@��m?؀>���0A��7�?kբ>�����p>t�~?��E�D�=��3��1q>#ꓽ��>���x�?%�`>����
u���-?WE�>^�Ƽ�T����z����>餟>j
+?� f>�s�>'$?�>��4�:�?��'>��+��ޤ>�cf?aY+?�%�?����H��f�?c!����3?�����>	����T'4>��}��꓿�_�!u�2�@���n?���?��RB>�����&�ٓ���-?�?_d�?�(�>�E�>�z?`�/>�64?EQx?1�>��?Al?�z�-8q�%�<�
���=��������@@?\�Ͼ.*���>�j���>��%�(�F�!�`�.�6��*�~�.���-���)����>@��'��Pn?J#0=1@'�����w��@�?�~���s�XB�>M��?�bZ?�8q��s?�=�>�������΋>孒�OJf��.�w�,�d4?μI�b�k�-+C��1?��3�]�+���=�r?�n��龫�[��0+�WV ��ٯ�a��&���dE?4r��:������창Էz�+�?�.?�h�<�;[>�%�>��?�����	>+��>;q�>���>Kb���&��������y?���?h?����ؽ�1�?f��+�?1醽��d?~�p>�?��<��@�m�}�
RN�oUÿ{��>v��S`S�����U?�z1�]�w�7?LL�>	E"?�8����D=e@?�?�/n?���DE�(�/�>[
������6b��ʜ��?�
�=Er�������퇾�A�>���=<Od�oϒ��԰�%c�>�ɖ?����6�
�q���
?�>��[��=L�����m?�y?@ws>V�޽9A�?)����?ջ4?�ݭ=S0������?�0?�Zȿ�u>$0�>X��Q�8�z1�Z5>��fu�yk�?�A
@���?~��wm�>�3Ͼ�*X?��=�����N?�^�2$X����y���;�C;�ZR@Ø�>��a�kQ=�3Y?�5@?|)�?��q�m�4?�/>��/?�I�E�G�p�k�I��|���1V��YZ�k~<��Fvp?�;?\=�>E�ܾ�]�?e�?�x^;Mi�=�GW>���>U�<?��>A�����? j�?듣>���y:Q=V�?�1>^�����>��`?��/���Z�s\����� d������N�=j[���e��e��c�=���>2me>��B�@c?j?�ν�����>�6?&a>�ΐ�m��n˾��>,�k>r�>��#?S�����0������ ?f9��F	?ŋ$?���=��݋���?	� �[�o���r>'��$��Pc���	2>�Q�>� ��鍾�}�=�'�?�Yq?w�?5.%?����ߗ�#w�v�,�R>��=3��s&>���?�	[?r">���=쟯��V�>�I?0iQ?kk?ު�>���g�"?+��?��¾N��>��L?���>@`�>ξ?<(?���=\��?�@�?>��ja�>3?L�<TC俯f�=��2@o��>�i�����>�a?!?��'�K���>8��>���=�{?��??wC<8��=HZž��Y�ɍm?�e=>H��>6bk���?]Q��z> �>��?�������?L~�?Ԙ>\f1��++>c%?\I�>������;ܾ4��>���=�� wཷ�8=W�����J�mǲ>u��?|н�i�L����>���?^z�> ��>�h.?4���N�Q����?�!�FX>���	�N��%	?	��</�?�#����t >��-��w����?פ?��t�$C��ÿ?+�A=��(�[���M��3���>sU� ���YY?�����ԭ쾊r�>K��>�~�??-@�?=B7?cfY�_��?��5>e��?����S]>m��G�V?��¾&q��_Dμ��¾dsl�Hdz��� O�>�t�l�>�2�?~�>�u�?��N��z*���Ͻ�?-�����Y�?Gt�=N��>]���\q^�r�	�7��<������?p������=ǃ���=����@?��<��=V�>]�0�M��Y�.?�.<�(���R�O��><�d=m��,˿E>�p��躾�k�~:�>X;�f	�;o~���?lO��:0>2� �����X?Y彨��L|�>9�T����꽸�ݝ�<��&Ԕ��ο�3���>��ľR_޾?Qu�G@	���u>���"̀�[QP�����ԩ���u �G+��� ���	��W�<�jv���X�z��>}��0'>U��?I\�>�
u�{ј>�H�?z[�EY�>3QP���?XI���?�[�>�m?��?��7>�Ͼ-Y��h.>���?���J�����>	>�}�<�,�����>�������]۪��6�?5�����hh��h�?� b��T��u%���?~�?wq��}�?�_M���&���>����_���y�/�����X��a)½�؃�XJ�?��k��;���2?��L�Jm�\��>��?C�?��?�X�?���>��/�6�?]g#?݊+>h�Y�
���-�� ���*��������C�z��=Vpu�����>{ӽmGﾻF�_�}?ȸc=��?qf��Xi`?��M>�i�1@t��=��׾:;�>��?y�>t2?�L�2�AU�/��Z�1�����B��mG>f۾�3����c��q�����o9r��/'�\���g;@��ĿeB>F�a?���?B��C_�?��X��|�?|C?�L�>Xn߽��?��?��S=1�����>��������*I���ｙ�U>�ý�� ��P??a�������1��^`��_��MMq�N�g���N=r�����9:�?�z�?m�a?r�?��?֜R�Ha�l��ފ?��Ѿ�·����U� .ʿ̊t�e?�p�������=�;]��" ?�>���@;�>�>�_�>V��>hd�Ug^>>�m¿��Ӿ�}�>`q�>;7㾽�?��6�C�W=@/!����?�x��ս�K����X>��+;ձ/?ޖ��ѧ�?�.�F����-%>Ҵr�x`>��<�y���i?�U[�|���s��p�>>�о���ꇿ�J?Z��<IV��>_!?:��>�f>Ͷ��1o�>��پ���x��<��z�>"%�=ӎ�>)�?o�L>~N(����E�>�4���=`l�>A�n?�ħ>.���i�?��?(���\�þWw�?�ʘ?���6�A)&��92�]���'?���>�b(?_�g�#��M��V{?0��*LV��R?��<?7#�>M�W>�|ý��?0LK>w�V?�>��z?0̫>�xt?�z�?u
���6�����4?y���z|ɿ԰"�OI�=�j�>,`&�j��?S�S?����ʙ?k��?:��XI��BK�>���?3�;���<�\i��uy�?)�ͼ�;���d�?�A�?hm����>'?3��>�>w?EJ �l�A?l��>��6��,�K�@?�V?�:�J[�?V���7�>@�9�>�b�?6Sv?a�=.��>_�>�(�= ��ǻo? �V>���>�(� R���ɾ��%�s%�HO�ۿE�=�C��'KL�l�ƿ���?�Ȣ���f�>�k�>��A� �?�:?^2�?+�3?�\?�C�=��x��Fl?T�?��˾쨿T��>5��=�R�������.������[e=j3��/�Ҿ���>���?�ɀ��o����r�*�?�X��i����׾��?.x�?�x����a���������r�"򏿬D�>�=4�3����l���'>:C6��㿽j��J�>ʚ��כ���q�>��D>8�-?̠?�iV?;�?.+�?4������>���=%Ώ������]�!>E>�05�\���5�=U�q��%�>B�	�/۸���i�c���dA�=�Ҿk(>u䲿t ��(�>��&��}+>T�.���?-����Ѿ�u�[�����X�sa#�걿>i���i?�9�nrz��>)?�߮���Z?�)v�E�w��a>-�@�;�J�i~�<8.S?���e�ӿ��c?�O��:�����\vM��;#?�;?I��kE�>�t�>�>���=�G��Y">R�w�M��>~{��>�H?��k5����>p�_>�M���I?��?��7�R�P���˾kֽ;{�? ��]/9�)�>f>�e)�+��V�X?,~�{�O>�?$��3��"Ym�ߙ�l������CA���1����׭��@ ?���	��<3��$��?��߿��W?	up����2�??�@?|�T?ʂ?�*?P)?��>���>��T��y�>@�b��]x��(׾����
s�G�>��N?�]0?�y�>y#�?� ��D(���e?�B*?�־��l��b?z��-
?�7�>e�X=�)?��>�'@�dx}>��>4�=������g��!Y>�nȾJ�>��̊<�\�>��=�s��[y�>��?��L>����/7��˳>�ξ�bؾ�ے���n=5�ɾ�����H��P���e��u~��Y;�s?#�5
���3ݾ�:>n��>�u?Q��I?Z��>Ї���=�a�o�>h��"Y>L��>��%���(?K��>���>p��?��i?�m�?B��?��[�h��>�0�>�AD�����}��b��ה�q(���1?0
�?���:��?0�??[?t3?F�=?�=?�;,?ǖ�?s�p?��?d/�>NPA��y)�Ѣ���~�E�^���ཆR9?P?��>�>���?��?���>Y�y?ZH|? �潘�?�ɾ>Ob7������N�=&�~���c��Y�����s�?���n���H����?�d������Ɂ���?n���f�?^��??�-��ÿĭ(?X��?R��'���j�?\��`�Z��}�?��?���> [<��?#m?��C��%#?	t��B�g?�'�=�H?y����� ?C��>���T=;���?�
��5>�Qw>f��?��u?�/�?�>�>f6�?*��>�3>;�D=k`����������������S?S��>��<?Q�!�t�??>;�=�p,��o>D�?����DAW=���e�Ph�w�i����B0=��?�ԋ��T�>2AZ?�`D?dɕ>���>k]V?Oy�?¡�?GZW?!�4?��?��>3�G� �]>+/�>Gf�?���3*='�6>4��?�P���?Ӆ-��F8>�;���R�̭��G����־�D����,�G;���x��g?��!�ꊾlb�>�'�>t���ݾ �$�j�V�u�>�/�[e�?���?UZ�;4
�?���>x���Ƽ�w}�?��1���?]0�>�a?�&,?��p��&�>�e��m�웿�/3�m�r�O[>�Wf��i>�!�>�F��AŽ>4�2?T�c>;�O?��f?�-�?�W?�7˾�ji����?s�p�-a�?5@ƾ��+?Y95?������.>vzt>�h�)�վm�ͽG�?��I?@R��]侩�<G��=`F�?�kT>�Yžb?��R?�y>Thؽ�C��f��&>@�3���>Mӝ��@������=��@��ſpWS=-fP?�9�>
���{?'��>J��>�/N�$Rv�B�9?�)
�,W �n�B�Io�<�l��5�_?[�/����?/�>��(��$���p��?q>+�?�fH? A�<Ld�?*4�>��:?�x��I��>`�����W?>���T�Dѓ���]���r����N�f>@��>5@;��M���W�>��>?��〿1��?�J���'?D[��e���֣��*0���>5�ٿwu�?�ા~��?¿[>�c־�L]?�ȇ?�<�o
�xH�?�Y#��N���X�y�������@>W{?S�4�n�p�Z���)ȳ�{t8�_�&��#>ѱK�@p�?�6?VG?!��>>?_��>D��?ڨh>Y���?�-@�1��f��@��>�h�?1��p����vD�@���w�����i@N<��0�5��F��>���K'� )?П�?0�a>P�8?^�@?�Z�<>��rY�>첊�x� ?���?J�Z�c�.��h)������%?�A�K��p�4���Q�b��>xse?�F3?<S?�?5�>���>iݵ���ǽ�l�>��B>,�ݽE֋=��ѽ킶��+ݿ�Z�1�����=F�/��@р�?�KS�16?X�n>��Y?�U����> ǝ�ԍ�?%tv?�橿���>�c=~����"�>#��>�9�XN#?A,�>@��=��>J� ?up?7?&S�>���?#]۽^]5>[?�>�l�>pv<-ۜ>l��{ 1���h�=ƾ�����Z>ڊ?C,�=7�Ŀ��?�!n?�ѿ�0F��PX>�(�? %����=i�>��?g�>ژ�?��0>�TI>���>C��?�l��.ȿc�?�}=⠞��W��}�?�8�>�/Ͻ��ﾚE���ZL�ը�� ��J9�Ȁ�>o����m�\�&��Ϩ?� ݼ�?d���<���$�=�ż6�=��=u[{�0��J��<�ۈ=�s����3�u�|�uK�>t<(��f��=2*@>�J�=Ǜ�>\�[=E�h��=�
�����kp>:?�>5�ýǲ��ǵ���� ����HT=W���*�{�ژ�>S�5=A�
���_=��p>������ý:	齭�>�n�>�&�>eu=��>&;1���>�=|<ǡ�I��<A�>Ȕ�<�3���w>��">��=y󾛦�7�����X��b'۾�ws�k�þ;��׭�����>�ڄ>��=i<����
>��>I�'?�Z�;���<��?���=f�>XG8>9ٺ>���>�T>�:�W%���Rǻ�s,=v��W���d:�D�T>�|C<���;�3|>)�=�>�*ܾ���=��=$=�,>%>���=N@�<O�<���=�?<~�>l�%?�H�>������b�=$T�>Q⳾�%+������'m�kʁ���h�P���m�3>20��>׽'پY5n��?Iլ>���>D��>�L-�t� <���U(�/�w=�h��Cƾ���=��>����9=�a>��(�/��>��=E>&�<���=#���}i�>0�<[����pr;��>�"�>�N>�ʵ==�>�'���ܽg�R������=�E>-�>��ν�gX=�5>�2<>�ub��GS=%�=#vF�>:޽.U������sB�N�A�<��Jb��k�q�C�������>h}L�%����m>������%����!>hC�>ʹ���&ҽ `<0&�_����=�<=��A>V����`�׾���2��(cӾ��C��������pdͽ�:{>�A>5�<�o=���>�,>��ֽ���Χ�=�
��_����>�>��>���>:�?��{�ɽ���,�}`�>U/J�K�4<�^��ט�>h�l=�P����<Z�>�
=c�0=k?�2Q>F.g�=�*>��>���	��=�"=j�?x=��r=i�=n�>>i�>�0>/��>�Ʈ>*S<��=�/c�`��>��^8�p�O�ʽ���>���:��Z�C,C<�`�>^�Q^�>B�>>[d?5~�����S�>Z�>�s��SX>�&�>A�j>e���_ṽ�!�����������:A
�����Ԋ>E�=ǳ�;����8޼���V?xl���ѝ�>�e`=�����F?�A����p�#W�=�#B�����2p�j(���m���\=տ���Ǿ^��(�����������L>β<��,?����M��<�>Ѧ�=~l���K~=~ia>���=\����ƾ�ž���OY>�����>I��>Bf��b�R�������:>	7�0ҽ	�,��->J�>�#>�)=^?Y>Ma	>/|G>_D�>$�>�a��`�=N߽����ƽB�@�u�a�㠢=`7������Պ��	��ћt>�=ٯ>W��>\�>'�:��x=Z�:>\�*=`p#���O�&�=��>��>J�Q>�s�>?�#��4�=��kO�=�d�<��<Hj�=X��=�8X=�WýfK#��g><�?b��>�e?���>��%=}?6=q �����=&"N<�d���=�z
>�(�<>=�༥Ѕ<	D?"��>3 ?@��>-�>S+��;� ���V>�fI=��;=�_O=�F=����^�4�=ɭ�>4ԭ>Y.D>�!�>8�˼��ϻ$�>Y��Y�g����֖�t���k�=hq���_���������&���^̾$�˾'��OW��h�Hپ�j��,2-���3���ş���>ƕ�������>V�+>�_;����n<�����?��ݽ,�g�>�u�Z����Eؽ.�=
<P<>1>����������������ҽ\�>m��PF<��E ׽_��X���>�=�v>��g��Ѷ�xa���ܾ�8�>k
=�W�=V�=d2n>מ�%L��,���c>�����g�!����)?$`�=��c>xL�>�C>2W������?<���=P�/������C�:�U>���ڬ-�����z?f�>G�|>��s>{X-=�枾]pj�Ym>,��=V:I>>j�=�;a><�mT<Mcg��>6>6��>ާ�>�J�>���>|��� ��e>?������@��=�-A�]�e�tt_���<:�W=�ɕ<53�EMξ�L�rľ�7>���&zf=[e���`E<��.���>[F��=�U��/�=!Q�=o�x��aS�����;��F�e��D>E-�� ht��>6�Nѻ= 
�>W��@�<<Se<s�<��> �>�?Z��>7l��,h��MN �����${��뛡�U���r����;>E�(=��#��!�>i��^��<�C}�5W8>P���p'X�Mݴ>(q���|����)�[>�}�Fk���/��> ���&����<�b�=o���	՚=1��;�k�>�n�'��;ܢ=�k�=�ŀ�,�=��<�^�=�L��^��: ���ʥ���r>$ɼ�u+?-�H>g����>��F>�Q5��v�>t(���_�>P;]>H���Z�ʽ�|�RԢ��ۓ����>�47�����<���=�}¼
IC�ی�= �>Q�;�Ɂ�w�b����@�~=��羛>>���>��l>_:*?�?\"�>Z?T��>Qd�>k�O?��>��>�1?�	�>H��>^�>�k�1z>%
>Y�P?'���\-�Xr�>�a�>�a�� '>��}>RZE>ἳ��M���0���HVȾ꺰�X��~�����,�ϚC=�= ���ʉ� ��=� >H�d��?�ԏ���e�~���M�>	n�M�>�T�=*���ےw���>ڟ�;p�)<v��=�R)=��~=� N�f����ｺ���Qʡ��Q=h�0�0P���9�=�����G�d���|�<^����R���Ͼ�r�>��%>�u.>#k>�}���>��;�Me�+�y>��L�|̊��R>(�M>� �=�����|�M����"����"���j���F �7���'��}	>u;̽�q��@.�0�>*{�=���8	��һP�4g8�a��e�n�%%�>[~�=_�h>kvþ��*>)I>�$?B칾�q=<�U>Ũ�>u�
��IK�*y=���T��>oAq=�)_=O�>_��=ax���;>O3�Z����똽�Ac=_��=����J�V�MT5=Zl��h��=-$���6?����.O�����>��&>E���=Ɩ=;ф=�d�+����	��/�����ҾS�x=��`��o??�	������G>��5<��Ǿ���=ܟ�=���������S�����������=�&2>�Q��_>FY>턙=� >���>���<�3>d$�=+	ؼ�{�>N�u>M.�>C��>�.�=�!�<�U־:��>D��=�Uj>��=>��Y>�2<�A�=Q,>��>:.�>K�>̊�>��>?[��6?�y�<qB����>�J$>0X��{���;W�=�C�=0��>,�4��#=�ih�O��=�,���E��w���K��0���X��G�=���=�>ֿ�+|>��>V|�=v� �h��=�՘������Ժ?(�=T���� =e2�=��9�4+]=�Nh=�^�=ɀ��*K��&��?�>�� ?{4�>���>W>?س>��J>���>�8���^��)�}p�>�?�YV�͌!�9��=p�8��R�e�𝉾��e>ጯ��[��V[��P��5�}�4�$���/��B0=����Ȧ��7���HD�n����7��n���Rf�����ĝ��->�B>ѭ���u�@�=�)�>96><!��Z��s�=?,*���ھ0ᅽع���*ƾ/)���zD���>�1��7�L;�[=yI	>f �t����8⽨�ܽ.�?��>x9?���>"P	?�ľ-^���c=�\�>&v��"�(<)r
���="c�=����_�9H~k��X����p��+R��c>��M��Į��ξ4�;�ɡ��,��~������>	���s9��瑆����_�U����~��*��Q�	� d���G��������@V���|׼<:m=�빳e�=,��;S!> ��=s	�==5�=i��<�S罔E���e=�f�=|i�=���=����.$�~0�f�Ž�pٽ�-��GB����=�ؽ�qʼ��@��7��U�3��D��̽U6R�O6>3�>�S}�WUc>�b>�����}d>�ѕ� S4=��=e;�=������>G�z;����";����=/"C�?�@>�O��a�<�/�N�bZ<��I�J��<H�<��ҽ���=�D�"�=ǤK>����$)��^�=�!��z>cV>˕�=�]�=$CE>���=�<Ϟ��N7��['=φ"���t�2����==gh�k>U�=�k=�pK�":�>�M˽��=ꆤ<n|޽���<�2�={4�'#>�$�=��;>��>E*�>�G�=� ս/,��w�5�=����޽�A��2;<�@���� ��jʽ�%S��ɨ�9���%�F��@�>�~>�y9<���=s,9=Q��=�
>�FʼF}>Gѣ�W���C���~;=���EAk>��f=�P����]��h(�0�q�>~�QJ�$�>�#�� iL�hۼ�ݽ9���T=+y�=�eb>cd>����N1=�%>2&Y<#>���=k�=f��=��5>�w�<FP�=i��=��B�&>��x<��;�����Rt?=Δ�2u=|M	��8����U� �|=�<㚝>Ю�=C���@�=����/C~��Ԛ=&�>��=$��U>�U���K��f<k�`=��(=�>v���7~L�t�0��Ӄ���_�:M��2/:��<9(��=�on=f�!>���<[�=�%�=��=�A>���=�B_="��<�$���vh>�e>n{�=�b�=cH >�^�[��<8@���_>u��˽�$���n�=G˽\�ȹ%m��ZM=���=���<ŦK>F� �T�N>u�<�TU>Ԕ=c��=�H<���=���<�w�=T�>9]�>��T����<�1�S$>j�d��փ�>����K=� �(�%>*MZ� ��R�~;)I���{�D>�/�k�>^HF=��i>���|2�=�+���ϲ�I����a=N�=,�h>����������M��JL��<�Z�6<Z��jY���\{�=�o�>��Q��
�=�7�=/�0��u�� :>�b�=<CD>�#>�d� �<�tC����=��żp�F���<����=:/��M�1=��n.=��ǽ[���*l���-������
>���<��:��Q�=k���5�=���=��,�=��Q=^�5���	�>����������?�=AŎ�7� >��<3��do����F��H�{���=��(=��;^SF���<.u>h�=�==F<>�cS>����ʖ<w����<o4��ؽ["�}���s߽� ��"�޽�W�=�/=bۙ=ˆ=e>��@=w尿W�ȼ��=�ؽ���5 ��d=z<Rť=�S�=��>U�1>���<Q���������e����@��
��=�A=1X>t>t=q��AG�=F�>R�<>�'>�>�P�< {̽����b�;�$����r����=D��:9��=M=7Ͻ����=��j>�i>v�>��t>РѼ�RU����yÖ<�X�<Vg�����9�{RC��Q��  =�ݘ=TO�=�>�
�=��=./�<�9�:ڕ�=�7f��l��Z�90�!��.���$Ľ�d��'	�����괽�rh�cU��EW������Fa%;܉�IP��n������<=6��Ͱ��2�f>ڛ�"N�<'����o��(R����O��P/>��C=d(@>��<���=d_B=���������w؏=ud>(硾��g�/��n��J�<�>��=3ռ��=�U�=v��j&<b���2����WH>ȏ�'m��.��2㽣1!����=�b���>.�曊�R�C=8s�������.�|@�=�x�5 �>��+�=���}X=��>:d>A��=m�=������=E�8�<=�L�=��u>�b��&�<�����->�W�=��w>׎>���=��̽٘�=�;U>Ԑ�<���=�՘=��>�j�=����U3=��=�]>�I^>T��=h�{>tj�=�c�=,'�=dM�=�o=�!>؄����*=�޽&�
=a�#=ź=�x�_�&�0���|���j=;m��V�<���=�����`=J��=�m=��=z!0=�ʵ��
�<������2��=d�=���=��)�n=&U�<��=�%�<*%->�.>n��=_��=��>n�|>�>��>S�e>��\>��B�(�B�۩S�;㽯bG�#iϽ���=��B����x������*�0�H���#��5Z���s��v=���<,E����=�W�Լ�EA�"��=I .�6S�<�����Y�<c�P>Y�<� ����> ҽ�#���>�U|>5tx�?�D=���=f?�mg.�3㜽H[��"�>k==���b��}�4�Ԫ�x:>"��=���>ط�=a��=��=�b�K�f@�=�=6�t>���Ӳs��I���B�eP=��!="L>Re��n�=n!�=�Q	=v���I!>�+��=��=�p�pN���p[��Ae>�/>�� >џ#>ڃh>�m�>m�>G�>��c>x�n>�wM>��=���>�
>��>eF >����;�W(>��[>�?f�+>0=�Z">��Ͻ�J=�W=� .>�ʽ�c޼ �ɽ�=��)����q��b��4׽�e;Z�B�xՅ���X��# >��<|'�;����L�]=P4
�������)>�k�;�ȼ=��$>���=�s�=vo>  > ��=
}�<<�����=!�+��1���x>��;S'.�y.��p�"Xg����D����1D���Z������ �y��}%�=�h���Ul�|H=����6f��4~<�G$�ꔂ=�����t=cJ��u���m>���<�i���z�V�P�k�9�.�"�-l3��$ʽ���]"�a�=�7��d��=�!U��=�<�P�=���=9y�<U��<nE��a���%1��$�;�c�J�=KH�n��=�=`����+�_W=�,�=.�T=���(��:�;I�M������j��&�
��S�/=��
��)�4v����ħ���D<����v�<�!�=(QS��|�|�1���d�f�>Bf�=[u�g�<q�=����$�D1,=	�@��52>�ɽ}�-�����Kà���v�#ٽ��=�=�NZ��k[=����N&ͽ0+�F�������rA(>�De�{�~x�Ne�~�=��	�0�V���	�b->=á�����=1LG�ȳM<�.��(����>�e�<0�=��
>��=�o���ۼ��>����=z�c��W=��U=���4���d5���<s�\>�>Xˑ>�3,>yv�=��=��&>�n�=K�=2Y>.X>/�!=X��%>�j=&�=>�7={���9�=����བྷ��=v$,<O=�=� =7�>�9&>h�O=���=���=��>~Ɵ<�|Y=�x-����=�9D�����X">hah���9���=esѽ���<IlF=܅���q>��=I >�4p>U=<�=�M%>7��=�}='�X��Y�=I��@`�<]fн\��<�W���e��D��=���x=�5)���>Q.�=ú�=lϽ���y=�y\�.�=����?�=���갽bD�<�����[��<1�̽v���-��R�����K��]�;L>T�=矼<!��=@�>}>|ş=�:�,>Wz�J>�:3w��)B&�󚲽_���g:��I=���)9��ø.��YJ=7�>&D>[P#�� =j�e��-q��K�>���>ь|>�F�>�2�>�̨<4͋>č�<�_^>̳;=�\��!�ڽ5�4>^�r�s��=CD�=�Խ��>�/%M���I��������d��XQ���=��ʽw��<6߽Uƨ=3Q�<zü�W�~q5�Og�<�~��E!��=�b�X����H#?;�%�a�?Y�?���?��q��S'�2(1��Ŀ>"�s?�<N?#���у>Js�?��A��b"=_g���hN �/��>a{U=<l+?���t�өx?�r˿Q�������|����9��w8�c��>4�>��Ҿ*��>���=x�>k-��N3?�1����\>�S-�Jړ��e�?�w��;�	{\>.��?t7m��FE�X�S?'�տ�혿�Q���q9���sl����q^��G��NI�qp���lھ&��+(߾4^���i�T�7�	>�G�'�����?�A?n�0�{��>ף�>ȟ�>���h��d�>�8�=/˳>8	T�.��?鑿j��>/¾V$��q�=]��<��`�$V<��O����>L�*Uo���l�G�8�>��?�7�?щ�?  �?{`v?ñJ?&wu�R�=�0J?as/�n���a4ľN ?ɍ�>�ZA=�5ؽ�q�� 8�=>�w�=�U��p�>�>�)ǽ�6+��i&���Ⱦ���>�*��֎��鉿*j��;���u�>|����`>�w����
>&d�z�޾�лb���/h���T���<ؿ�?8C�A��>_?�ޖ?�:>� '�s�)=�%�?�I>��
?O����3�q�W���?���N\���=�5*?�f?s� ?-��r�)?��T�g`�b㏿���&��/ž�,��a��=3"��������#��=��9?T6�>*�=r	׽���>��>�ti>ċd?��o?@�>l;Q�`?�>�F��c?���>1�'��P��P�>��ʥѾOA���]>tko>��>7g�>55?}��5���!�ԾD�6�����]�`�[\b�Ä?��>� ?�8�>o�<�"�?n3�<'܍?�)=O���/�=�����>�^>ߦ����ʾ� $?���Tf�=)��>�Q�By"?���}?���_C�=����-cF>3���J�o�wG��cŧ?�B�Ah?��|?u^�?��<�����ξ�=��v?U$�2D��B�+?ܪ�?:{�<3�UǊ�N�M?	��>@���o>8#>�3�؂?gE>.�;���9=��>��>!?�<�?��>��_?���/WG?Y1��g�M����v��`�`>$��>��3>��>��/?�1���?��#:>���> o0>��A>��>\Ϊ?'��?�Z?��>o�??��>#.m<_r�?�K��ݽ�=A.��
��UѿN��_-������W�>r�C?x�v?�1����<���>2��w������M?g@̾��6=Z.��1>�%��K���Ѽо��=׉>ۿ;��I�=gfo��������>��>��7���̿�d>���<�==�9-�ln?qr6?2�E?���?X�n?��rb?W^?m6�?ɥ���H�>�E��>��S�W�ҾA�������;?����?�P�����>{<?�*��<����z>�N< þ�����=��پWu�?�)�1C������Tiq>�1����==��>�`��͎4>5�(�6)���uؽ S>ԝA?�MO>���>�|���`��s��~��?��D��Q�?o�n?}�@;��=`$���/��Z[?�<=$�u?x8�>Vֱ=E�=����D�3>�Rj?�x?�����_1����@~�H�葾�S)��
�>R�>�� �]>[!��L@>�J3��V���+|������-?��d�k_l��3>�� =j�վ��%"�����=�罿I���$F�����JnL�X��>��7=���������ސ;�7�Y[־}�>䤿�6L>G锾��>���>=��>8�=>��?q���?^��?JƇ?���>Q@�>�{3>1�A�S����K�`�!���!�j3�?��g?ܦ?K�<��Ž�Sc?F.��Δ���y�>[L�?T��>a�?�a�=��پծ?U

���k�%ӏ��>r�=�DG��E���B��N;���Ŏ���S��V�S֒�W�=63�<6�|�TK�`������,=��ܾ�=|ג��b�k�o���<���P%���|��:?؟غ��:�$V��Od�� �4�?M�e?�3���[d?��?b��=����e<_���r��ȑ�>�I���?��q=������#�T��3��=���>P�=��>�׽�է�b����Q?�����Z��AؾmdT�������
@?0��>C�T?�.?Su�?� Խc�l��
^�JS{?�68>}d��!�\�'U�>�Q����> �x?n�^�[Nl���>�,�=�:P>uRB>���>���>��H�w8��;�?e�=I}$?��%?V->�}����^��E5���	�y�7�$�F��N���i���n}����2U��96��eO>m��>tl<!
����K>��
?�M?���>�,���0"�S֖?��'�K���ٍ�S8�?*��=t�S?A?�?�^�?�
���,w?M��?}��;�=��?{��?���>W<V?�?J=?�^x>���=Of�>�K�?������V���?�ڴ>*��>����C�>!�Q?+!�?���>=W�?_�Ω��#H���T��Y�*H7�i��?��Y?��?���<SP>���>�1���K��ۘ�?ö��Hɍ?�4-�]��>?}߾YdU?<#X��x�>�H�;�t>4�T?5��?�?���>)>�>�'?�-?��*?
�?Shb=��?ȃL?%��?����Yq]?p��?���̿�R���m?�F`Z��о�t�?���>�����K��_ї>�>j!W�bCɾ��d���=(�J�$M>d>��">��6k��z�=qO�>oq$�bT����������b?��4?�
:?�
I����>�/D��i�>�P,��2�>��ľ��V>��}�����D��6+��\`�Z�+?�::�>m�=�[?��>�����%���>��>��T�!�?�/?)t�>tU�?��?7�=���?C�#?.8�|a>}f>-ۄ=��>X�>��?1���9�`2�>x;
>nG5?��x>Y��>'�?j9�>��ۊ?�w�?�A�>T^>�T��>qL�>Ϛɾ󇵾�L���>�L�>?�1��g��3K6>��W?�4Ǽ�邾4s���i>A����\��ц=�E?shl>�d��C��>�1?�����:=�B���s�o�]�������ūO��)3?Z���U?��?()�?�"��8���:���>zw$���8?'��?�-���C%�ʬQ�r$?����x?�G>�y>�n�=B>龅4A�;;���b�R�2��z�>�~6?Je��b��B%�=��8�M&"��;:լ>���=��'�?�R��T��ZM
?{脿��=�;��C<ᘾ}�R���@?7칾���<L�:�^B?�վ%�e��j˽�E���C��*��h��8�F?�X�?�*�{�R?Q5>02\���pHf?�c	�$�v����>RL
�_.�߭-?E�?��n?]�/>�R�>=�-<p��>�?LX�?V���z}�=���g�@�+���:L>>���K��2���'�>l�?��Y?j_̼1�/?pΙ?Q�D>P�e���<�[R?/�>gr?F�?�=>��?8�?y�m?6ŋ?0tI?���>�|>J��>�ǘ>>K�@T�>H��>E�Ӿ��:?�FK?&.+?�A
?|�?�*�>�q?�y�?Nq??k��Ȅ&��;Q���J�[n�=#�>=�c?�;�>��?��csʾd�����>?D|�٘W����a�%sY?>��l=�������>x���I��Sq�=����R��a�>j����^���>�5񾵼?4C������b��'r�k(��4?����y#�ǈ���*?)���Nˋ�������Ҿ	�M�z�a?�}Ծ�G?�����`��,G?ԝ�>	����>z?�C�>��?�<�?#j�?nOT?u�u?ŕ	<�IV?~9�g�?�gN>R��KT��.�?����B>ߩ�=d6�8i3���1��Z>�����s���C!�a>�=�H���R���c���þл)?���]��>ܛ������R���������G�>񐂿nh>:�x�|��&�>�#��I�+>�Ԟ=��>�'־�	��e
?�C{?�?E��>��?�?�&?%�?k�?�@�?��>>��OK> �d=Y�=s
�>��=��L>��?6W�>�����5���7=?�G
���A�x'[���>��>�D>)|D?�G�>K��>�d����v�Ƞ������j]��Ns�b�B>Fp�����~�A>[�ǽ.����̰��I}>;��	�N�Ӽ���k�}�>2�Q��A㾗��>�B7>I�M�ߡ=��=�(�>9�n�x�U�J0� pȾ�)�>�"��>X>��,?�ܗ�<���7�Ҿ1��>��r�ξ�n�:��=l%���
���m��}>�&���6�����{T�>n��>w�}>*��>��)?<Pƽ{9�x;�=CR?���>��,?�Z!?@�1�¹6�[jd��zJ?t�����U�6b@>M��j�>B�����=�>e��>�@V��⌴<�mA>�H_�y��ϐ��u�
?��?+�?Er�>Г�����>FcȽ����Qi�����M>�DN�U�e���.?f��?��a�e�u=:2=n��>�#���{y?���X<l(>�/�>��%?��˽�;?tվ����܌���y=�E>�����wm>@"���=��<�s�A�H?��1?E��>"$���꥾�^���0>�Q1�nX�7���o�;W�>��ʾ$ž-�R�Y'ξO���f�_,�>�>-�{;�>��#?
��<��>k.�UIP���j��TO>�A��ʡ��@>���>��˾#'���˾9�����dg��O��=��U$�V�>e�D?h#2����"m�=��w�U �/w������3>� i���?�B>����e	?/��>-�L=x��gJ��Ow�>kp��b�Y�4?�Ũ>�����>}�Z>�𶾵���?e?����g���N�>J��>cL�=��d>�/�>��>?��˾��=�̓=�(?�{*>�Y�>&6ؾ��L>)uH�����(>���=��;O|?��{#d>"�>6������_�D�5>C�?4�?�?mn�<]�=�^(=�C?��޽�Vc>�1b?�u
?�h�ĎA>�#��νK(}��G����+*��>��,��>�F ?���>���nM�>�8>���Xs���_t�#��>�V/?�٢>��]>O�`�>F>W�ƾ;�����>{�S>|���g������+��O7> �����>��g?A�Ľ[�<T-'�r?�P�>���L:�ǒ�=�<?ҲP?W�q��LȾayI>���>$굼��"��A;?¢>��	�k�3��[5?>�������Y���z>)ʇ��[���O�>|-�>��=�U-?�L,?�ε>��0?g>�:ľ�o>�ը>�վ/��Ԉ����>NeF�u�4>�%���X~�=��.=F�D�"7�=ϥ�=�	�ٯA�$3�=�q��ܺ��+�b���$3?�m5�T6���/ɽ�
>$%+>�-�u�ƾ�؆;��=x���7v+�-c
��^?�w�����ei?)��>KC>Et�>��@?@>�=)^�?f�����(?��h>�V�X���ƾW�?��=�h�>.��>��N?�P?���>0򽪏�s�>Q���h�=cf="*�>!�?��?>/:W=(�0��8>�T?�,1?Hpq>EUO>��=|�����J��(*�_��U��>�
D���/�զ>���C=<�?�����}9��e? �#=\�d�S���O�PlվK��pP�AN���o�>���m�v��%J��b>��>�^�. � �_>�$!?��>���������v���,��5����$�6"V��^��s���A#�Oe��%-q���?Gd��b�?��j�:�+>n�V?�G̽v2�=#�>?2�����>6پ^�7��ƾP�־�	�=Ձ�>����5i�� y�>��������4Ľ�6��VH�o=��a/�!�`?��M���ᑾ�ˮ�Fɾ�D���'�1�3��?�<��=v@��澽83����k��t���{�G�#�Q�T>vr>=S���}�ݾ�ǚ�)�z��4�-���t���q��3�8	�"��/��(k��N��X
�3�O���?p��3B?�<�@������!��a�j����=���>)B�>=�뽚"��ؼ�w��,O�(��%�����;�0?�>Jw?��ν��?ϓ2?p�>ź��U*>��?v+�>�;�����q���_��>2�V��-*>ˀ�>��=%[?�棽�����b>Ŀ�>}u�>�?$�??�D�[����j�����ž��r���Ծ̀H�z�V�8#U�t��-�E��>?P� >U;^�M�i�4�ۮ�!N?>	�ξ<�a����;��>�Ӿ��@��U�=���>N�*���=�Z����>O�<p%ƽ�>G,�?U�7>4g�?]R>�t2�@.�F�>_L�?��?+P��G��I�����=Iq�>�پiK�>�B˾.`����׽q	l���I=g�Y���1����>a�7���d��-1��+���`L?�}\?i#̽1�D?�ȭ>�S�>c��;�D�>�3=[�>��,��Ҭ=@6_?ؾ/01?���<�e	=~�x>��>�%��p�>�� ?#F�>/���V&M?ڏL?���>`>u�>���>Axy>ڑ�=Fm־�9 ��=4�`?O]�,kI�즼�]?�[���]<b��=<��;9J?�f���C>fP��	1���$��"�m���]��5�>:�>�O���X�*�=���<�����ž�RN���+��l�>5&��� �2/�>�r3��h���m߾	��>(��)E?Y��>�12>��?g��^r�=��C�	������I���q=)nU?��>У:���ƾ�-�>+k�y-�-T���7?^��>�] > Xn��2����п�5�> ��>���I�>�~�7���6�iN�=0	7?fp���>�^�=пz��/v�+�ϯ�|?��Z�������;��>3�<+�>P��q}ڽF{����>]Mh>U�:>3e=NB�E
��>)d?2@��?���;��>r&�I��v�>m˜=��C�� ���ǽΥ�=��q��4�>��>��H�S����Y�����?ӷs> ����s�>P�˾>��D���=��'?Z�U<�� ?M�?%�~��^?.)?�V�>���[?u˾?��>|J{>�4>ll�>�a�>�RH>�d'?�e���(ݾ4��=�L?�Ƚӱ&?�1?�Z�=ih>��J�>j�;��z��QӼ>�H?�B�>��F���C���='0>h�[�a��>�!��8?���k�)�>�,?S1̾A.=<Q袾"�վ���>E
?��Ѿ��S�{��>���>�?*�>F�ˑ��T?�u�9�`b�qi�|��>��n?�����ͼ��,��A�>���1��ף�>Eі=����0ܾi�5>D���u�<�n2��{2>�?t��>̀%�@|�>ֺ=MV��֓D�'��>�=?qJ#��^����>�9�?肈>�t�M8?�֮>��<�m	��@?��?�d�=i�f�����ct?l�x>G��=B��>��<�F>�v�>��f& ��Z����CL�=�־X�>�о�/T������� ���2��!Z�=�ؾJ6���Ua����>����t�����oMj��j���o��%��=>���5�����?������]	e�
f"�����H�R�?�O�Q'����Y���?>l�>)�>�n]?䊱=b��>r���܋�>+�?bY̼:4)�C�s�N�������U����.�~��>�z$����=��=Ya�=�.��3��>�R�ó���ͽ>��>"���-���͍?�)�>�9������>3�>yl��V���x>D7?3$Y?W6ƾ��Q>D�������2R���V=AdT���R�!,�.V������_?��n��1�?N͌>p ���E�<��?�ƾ���r��X��@L@�� �귇��ؽ����˗�2��y½��>��.�."Z�PC?*��@����)�?��>�q��a��O�>�;?�s�=�Y>�ׁ=!x�>���I���������W���ŀ�o��C�V>�v=�x���j/�j�$>�-�>�m	>.�+���M>6.?L�(��'�;`?&k�>�� ?�]@�=��MP>�o�?tw?2���\O?%�|><�l?H>佫!>��>G&�>��-�����q�ؿM����p��-Ⴟ�?�����s6ڿa���|�0?�= @yr�=1�]<ل1?R?���=ͭS�y��>p�X?�1�9z��Pnn�׬������'�Wu1���>��@>*�N��<�&d?>�?Ϳ���v�-����þ���?�ol>��i�z@�>�P�?���?'��?�G�?�P�>XK�<��5>Y;>�2>8?���#��}�?�RN��f2?���>M�^>"z��v�ݼ��#=��=C;�>�ӟ>�d?��>ǖ?v�q�@&��U�[�PGQ��v�چ��nŒ����?�3>��������x�?��Z?�L�?A C>��f������7?RY���?t��?�K����- I<Vއ�T�J�b>����|��S"�5��>����-l&?�x?���gMK?Tlq�%�>�9>v�T?��?E�T?c��?M	d���?e��?�\�>��A�<��I4����0jQ>		-���?:�?k^_?o)+>Ygu�N�?��j>��4?�� ��.�>D�?�=R>�˦>�V?U�!�t�%?���?2�w?��l�ȯ�����=�ػ���.��p=S��=���>|
�A�Ӿ3�<���3?G.��p��?ͻ?.�?g拾09?96?P?���>�0�>s5T>��9=��=�Z�=�K�=Ks/?��T�Y��>��ɾ�d$��2ȿ���>��r���F��5G���%��w��+��?��?~���X��L!�yf�?�B�c���v>�٫?��?x��?��?��?�(?�$�>��?�EO?��6>���Q�پB�a?��g>�^���ؿ��M��gڳ��B��	P>%o?7�>%C�?_��>@�?�F���+�?
�&?;%�?3�S�T$����C?X��=2N���q�'��&��=������ܲ�2�8���a�.R�>�>-�; �>���=+;�=�-�?��ȾV��>��l>���=��?[�@$�(?+����>���xt=~G��A(f>t'j�{�9�h����	��S��i䦿��
���U?�m�����>����H>>�B��>^��?��6�**G���q?1������;+��E�>�?�����ʾXjc?��?q��>�2�������]g>.>&�)����(g��` ?-��t�?ʢ>��?T��?1�?�!�?N���Q�0���ƾ���> Ŋ>AT��^�?0�?7��KZC�%��>��@?���>u��?2P��@_>� �>JՆ�)�c�]�����o�^��D��oѾ7h�?b�0?HΆ��ĽIg#��U���p����~���2<���<�}����f?�w��2?������m�O�1�ո�>��Ӿs?���d�V�{��"�>(Ņ?��6�Y S�:8��c?B��<w�E?���+9�:�������8�>������пi���=��?[��=:m�>5G�>���?"��>�o$?8�=�V?A&�>�d�>�2�>�������B?.ґ�9W�>%���QZE�eQ��|}���Ȍ��x>�q����D�*�?ߟE�Ey��'�xs?H-$�b�ҿ� =���qh�?D⢾	��>�X�?Cnþ�25�Z��<���?��+@=�"�l��>r�B?zJ���?�L_?�l�>���=�/>$�S�`d=��޽P���,�y�}>��$���x��Jf?��r>G|
>��>&�?�ھ��'��Z�>�w��`�?1R!>���^���;��g�\2ž�v���<�>��ɿ�	J���L��\�W@>u�?���O�&���w?��?qBS>�<蚂;�i�� �?�����=����$���5�wE@?dJ�S����~W?L���Ƶ>���>$�� ��@�?:�����?��>������#���0?::�?\�H<TL?�؁=���OU�>U��?Sƿ?s]�>=	�?fΡ?7�5?i*�?Y�U?H�?S����?'"��'�5��p�=q���:���B���>(��>C��pc'?��?�%�>nd�����?�̬>n�ؽ)]�?�k!?z�����="!�>x�|?��=T�>�m���W�����j��GwZ�T�>q�5?��?c�?��>.�<��>�nK?�s�׎->t;��t�ؿ�R=x����?o�/��4�>�z<?�M�?�=T�H?7?>�=N���<��֥>�#=�\?í?KS�>�E�=��2ś?uV>�Y5��B�vE?:�>��< ��>���?��[>=�@&E�?�����7.���@��?���?�D����)�h �>�c�����a�?DG���'����>hd2>L���m�T?G�A>�8!?�����1?j�����?�Ҿg�R?��P����#��USh��f�?�� ���?�E��[.�>6�>ru�����>9g>�ML?Cm߾"��
=�S3���F���6�٣:>���p���@>�#�y�> �y>@��>��?~w�>�����/=���<ǊD?򀾚?/���@ʩz?��?) ����?���>�֋?8�Y�V��>C�?�I?���{����j�5�=��R>�ܧ>o�Z������i�?���?�W�>*e�=�I�>��?�k>�`r>�R>�[i����=&�>jɠ����>r�J?�b?����6\�?Z^��[mR?%��<�⌚>�xO?m��U?3a@=;�#�tR��/i�K�l������l�C�v�����*O7�8��?�x���ᶾgP����W? �>%j#?G8?�{�>��>�[�?�@�+o=���?^���	X���̾*�>'�Y�h1�����<�>�R׾��ѽAS�=t5>X8��{��;،��ξeq?��z�"?11?��>�;ܽ�j[>��B���1��$�@���d?�-��{��>���!�:@�4?"Mg?� 	���=#c�#��=�Z꿄�nC��G��6_>�2S?᳭?��Կم��-�����mF⾹�>5i�?�Mq�ȝ;����>nv�����,�� @N=j�?�$�:�w?�{9�B(&?({�=�9?l0�:yؾ!p����������.þ�n��/>"�=�x?ue�?���=`|J��$��k���?��=�d�^1��ޟ��/���|�ش�����>����a|�>�@�?,4=>=+��&U�>3b??%쭿`�5?`����8�I��?~.�?� �?^�e����>Y����
�<�V�Q���^x'���.?��?����a� ���1�"�h�Y��)��+<�??a�?�+;?��?�_D?1;h�8�7?��Y?Ӿ=,D���m?6I�(��>򤋿5���~7D�Å��ヿU�g����_c�[���%�>'/�?t~>G�?���"�>�In?�#?��b��U2=�>lFn?Nx9����������WL?���>є��;��C��>�"l���1?��^h���r�=�	����N?�o�=����v�|>f#�<4�j�l ?�C.>}b��V$N�9!��
�Ͽu~����?�͟?&R`<u���gk=_���?XVx�c��>�!�?ڣ�?5�S��)�?q���3��>�L>
�>A�M?�b�z�*�o�
���>w���%j���=K/�?�K?�(K��l��B#�?�(�>�б���Y��T(?*��c ������1���>��<��+N�ϸ�о�\��J��=� l?6���(�8�p?�K�>t�տX�y��RM���&?��?a�qN�?0E�>2>鵌>��=�����≿�����kb�L8�?���
w >�̿�a'��D��AV?��ֿ"�>��2���?J��>^��>@�#���&@0�	@�*�?*;X�(��^��>����1��l�d̢='�>�W�����>����H��oY���,?�B<�gY�>g}0?M8)?*�t��ֽ	?!7�>�^��B]?]/G?�d@
�y?�ײ?EU?L�޾�T��%�ͽwe�W������>8J�>>=��;�о��ھR��ӿ�V?��n��?�:?Y/����?$7�>Ek�?��
��W�?�_ÿ
�?�c��b	��	�>]�>Qr�>�櫾�G�?�	?ZS�>�A�=k�1?��(����>��>tVm>�s>~�>�M��[}��߁N�O�?M��=)�C?��\�>���ws@`Bg�B����@�S]??�-�[+��;羑*�>?�ٰ���R��D;��}�>ܑ=7�����>��>gF?�>)���?;�y��]"?��>x),��D���h���3��߾h�5?
�c?�W#?E��?��!��&F���������=}]:�.����þ�Z���Ľ��房�?bH�>�\�X��s���>��!>}	���_2�2���z��X�A��M��`�%?�<)���U�g"d�y�P> ���U0>��>�<��9�?{��/��(����>�)�㿦?Nֿ�/m?U�w��-�>�|?�=�?n���$��? }���I�>�:]��s?J�>�R��J��=l�����e�1���j��g������L?Ve?H�>nJ�J;����>׭
?l���s�=D�>oo�u�?h?��ʾ���~�?��s�?�w�?�~�?�>�?O�>�����U0(��?D��=��G?��>�^u?���?L.��~?o��>σG���w�~n���鉿f�N��s�R��'�>��,���S�M=���@�R?�-"@��t�'��?����g��=�Y?���=�:�>��W?ѧ~>s(�/�޾�o��`�=�]-�*����*�^��=�����_� >>G��>�Wi=����a�%?7�羰�T���-?�>OB(��K�w�W���Z�������5�ǅ��1�?D�>&�Ǿs?���>�	?2�'�O̗�L�{>�;��[����??�w�>;�@��߾ۘ�������5;���?�ܮ? f�?F@�>��K?�A��
D�>3�>  ?5^�?1i�;� n���@?3��a{r��/�hU۾�a�>M��=q8��J�R?��>Òe=�v�N܉>�߬��cy�� ��%'��o����/;G�t�|U�?������>�꿆��=>ׇ��/�� 6ݾ.�X;�"ؽ2ʱ>qI��~��>5��>��"��%����?�]���i�>����<�(?���>b�`?_^��~��==�T�=N0%?3?�O编)%?�;0?(w�>�A��Up�?��(?"[.��F��o^�/l޾���y)>H�
?�=���u��O��s�;��o?�|�?�`?�C�?"v�>jM�<J̿:��u���l^Y��t׾"����?#�ƽX=�3��οf���ZN?�4Y?�ɼU踿J9|�$�>�x�?�#�>�<?�e��lI>��?w�^?��.��a�������?�e��(�q��=��?H��?{<�?}���F�L�/�A�>đ�?1z�=Ф>�mj?��ſ��ÿ!�&�5>��\?Fd[�_$?g�ǿ�$D���=J������5Fi?���rM�?�T�x�����4�&@V=v? ���2>�䲾Ϸ��6��-۾q��>��S?��?��?u?�6?7>�l5��6���������?��7?��?������g?[<�>ܵ�?�J��`_z��(���N@�����*�?�2�?T>��U�R#u�,
I�[���/�_d��M��<z��{$?�uV��v�{��?=t�?���?D8>��G@�����������?A:�?-�?��?�C7���c���X��������?WP�?�$�jd>���O">)�.�Cݏ=2�T���B?�gv?�r�?��>������A�[��.8>����c��k��־X��KϤ�u+��n6�y����ڿ�A��'g潤�^�F�g��R>j�t�q^�>2.��{<�m�h)8>I��>��>ˑ=��Y��;r˿^��<�������=W�?���>�ش��?���>b��> [:?<�r��s?�2�ԓ��w��F��">O��=լ�>$J>��O>�C���(@��?�0?{'�>�>���͈�\K�?ܞ%?VRؾZh?4u0��t=�3j>�%���F?[�?ȉ ?��?Փ$���@:��?��>��?}MB?��=�e6?bp�?X=@9X=?	xh?�����k�("?d�?��>&;@>Iļ?���8�?	�V?o�k�6ٿ�^9>1g?t��?L��?�9:>r��~ۿ���27?��?w���H�hV"��!f?̜��B������k>s�S>2�1?�y���o���S���L?�1���X��7>���?+<>���$�Q��?�m�Mr��437���?����=��?|;$@�7�<���_��?���>�#?=w,���}�?'�?"q�?��q���C�e���1��o��?��[?j� @x�F��Y��.�S�%�f���=�D�?���?�h~?%,F?�&9�U�'��E�=�T���@��!?� =����q�>�{�>��P?���u?� �>g1M?g���'�$�J�s?�	�Q��!w?�9?uv/>n��?���>5(?s��?���=�?eG?�ފ?K�a?��h�ڻE=��>?�@?�km���j>>��?4�?�)��9X>�kýI�'?ƥ��%}����#?;�>xꅿ�Iο��(��+�J�=��>L�S?�5+�j�����>.��<�>�Z���z|?#�>����<���嚾e�&�Y��?x�$�Y�?��-:��,�y֯���>:@L��M?�;�i�X?d���@�d>���!���飿�
�ԝ���x��E�ҽ8�>#��>FQK?Xx�<�!�^�ȿ ���V���?��>
�5>e}�?�餽wU?h��ui��Y��߽=~��0-9�U7�=t��?����_QĿ�<l�����UV >`{���2⿟����?�?c�!����?��>Ps��K�� �x?��W?(y?tJ/?q	�?�P!@��?D���Ͽ��?����?��Ѿ��L��(��,˳=�p�? ���%�?a>��H�>�;ǿ�B?6��>2��>%���<Qܿ��\���y?q��>�z���BRT�F��ETv?�+�>/B�=R���QW?��G�97>ޯ�o��?�u�?-�ξ��6�c�v?��?�Yƿ��P���E�>^�E?|$K>[ �>&7����寿���<f�?E[���l�����ү�����&l�����u��!?�Z�t-߾�_��W����?�]?O�|?����~�=NqN�gMh=���>����B�?a%��߈j�T)0�o`��*ɾX\>?y?��ؽ�����sx�$���g=l�F�?b�r?Pk�?��@�8ؾ�2��0�ʽ3�D�	��?���?I�@���?OH?W=վ'�]���B��?ގ��J55?���!�E?�"˿�Ϻ�
�:�Dx���п�8X>�c?� ��>А�>��d?:�>f�h?�:?��>��?���Q*?�v?���>m�?۝k?�^�����{�{����=�:?6`k?�N1?&���R�>�z�=-��?�K�>��>��?��>��?�1_?i�}��E9?f�>蟐����r����������*M�>cs���>�>����>��?�@��A�>���?� �?	:�<�n?�M�?bkF���޽��ξ�W?�ᒾV�ȿ�
�>p�%�ţG����*׾>G�>���><>�=2#?���>4"�=�5?�?���?�*?��0?���=S侱E�0?,E�F�1�BK�<TwU��~��UJ?��?B��>/1?l�P���?|`���?g(��	��>r�?�X�?�S?ny0<�(0�$?�.~N���&=T��>�a6�R���@!+}?� ߾V��?�6�?��:?I��=�����K��{>��?:ft>��=���?�V�j���O+�^�.?��2��@��8����G�$��?v�'����'Ǵ�7v�0�?��
<��?��V���>nf޽Gk5?L׈=�E�z��M>�?Z�Z?^g�=@*�=ϫ>&o�>3����(�����2̿�?!t>�	?�C��Q�޾ԡ
��q�x�6�r{>;�>�*?���R��<P�ۼ�>���\�:�4�����>~Қ>�n�>r��>���?l�<<�i�)���ے;xD�>\A=?�|C>�Ұ����?؟�>��\; �fe(>(����$��f������4����)��1�+?i?��C?=z�Ɏ^�<��y���g�m�F>▶�e	?��>���;�I_?��*?Gw1>o|̿CTR�s��>|��<��(Ƒ��:7>^K̼ʜ���(��:>��>~��%��>g*?���j:#��������ztc�|i?�7D�|<�� ?[6�?�{�?.�U?��B=2ƾ%��<G_��`��>䋾յ��*�R�����ɿ"<��^q�=�Ͷ��ү��{�y��<X�2?H��>'`�>e=���>uC��B��a{����=Cσ��c�����=���>6�%��A��19�Uk}����?���.��ʚ��k���q?JG?*��?�P>aw�>'��=_�d?/�ѽ6jl�:�ӿ��˿�N�>~"J��j�}�?�%t��kF?3�k����:� �>�2>�?��Ó>��u���E?�Mn�����ӿ���\��ڜy?�l?T��M�þ �.<�|�<�)�a#$��c�<$N?�?U��"7�h;=ݨ�>-F�[M��?�>R����6�>�;?g�?�ܾG2 >� w��V�����C���V�<�}���*�	s7?��?���>|�I��[�#g$��í���"Cվ��?��}�c�E=6f7�̱ �P��=2�c>�_׾��>�X2?l��t�=�����[��>�_���>��པ�?��$�$�1����IU?�����=���>rw$?i���_�]�����GQ?�l?�l��g,?��?��,?�?
$�>��.?��Կ`��:fH�_�>�"2����tP�=�x0?��xn����a�܎>��4�b�K?��x?��>��7�k�>���>�B�?�9x���m>P���l�?j�������֦�O�]?��o屿E�]�핉��ʾL9?��>�~W?Ӿ4�����q#�H���Tas���0��Y<k��>�?���>p�>3ǲ�R�>��5�J�]v¾W�[����=rh�"� �G���Hþf�r���{�/�r�>Iq�?͌=�I>E��>90�>�U���9u��Hc�'e佅�E?[�;�I5�>}�>I�?������u>)�5>�,??4P���?��p9���?���>�v�°��h�>�i%?u��^�/��I/?e.�?j�~?C�)?ķm?���1p���h���q>�����=l��=��?�[O���w�4�G�W�`>���H>Q>��>W �>�̑�,�ҽ������>���=�����C>%A�>%+?ce��5�>zi*>Aq��"�y�a�?C�>�6?'\�>�8�?<�����?��;>��:"�a��l?�$�?Ѥ�>�'?����M �3�/?�V���z:?K��>��7?��>�����>�qh>�� ��-�>?��>�\�>:�%?JD�>m���{�ܙ�>f�ž�|O����ҽ�y�=�����<����|�>�G>-]=�q>[-�?�i?J�ʾ�|>�I���O&��6�(�=�Ž��6>��V��P�<�X�;E�\*���-Q�h���A�S��q�����>��p�>p�>5&?��~=↾�"�S��>Z�e?Dr>�4 >Z%/����>�J+=3������'z>��$>om�=��K�X�[�;�?v2:?ٻ%�q������-\��?�[�?ܫ���U�:�xW�\�������7,>�@��^<�p0>��Z?�Kž�ࡾk����i"��??2�/���;,,�>�˄>�!�)(�)�غ�T�,���{\+���̽Y��>��۽�L����؆�> �<g-&�8o�>��w>DM�� ��׾�Y�=�0����ؽ���q�>�w��X-=�E[�8��!ã��q޾���)9?-�>�����؂��ȾW�'h�[ld=���>9"���8?У@?%g��:(?y/��~��������>3��<��H<L�=���J��>ˬ�<E~�4)���&Z����5Ͼ,q��o?Xe�>� ?+��>����>*�u55>�+�<Ĳ�>�о�?�`?��?�ci�oL����E>�F�>�ɂ���<��H?0v�>��?���=+OQ���ؾ3e
?�/I?��Q?��2?�򣿔\����e�?��)>b��[Ǡ��	b>Q&�>�33��~S�6.���)?|ʓ<5��]b��'Cھf����l?������>?� >�~Ը���p��=�>��>I���4��
�?MBr>~��?12t?��4���c�!�]�Ɗ�K��P(־1I��bl	?V��>m������m����,�bV?�\?�ـ>��=i.p>��?M�컒?v>s@d���>,0,?�T?�2���h뾬�'�?�}O>?u�>NN/����N��>)!�>8u�>z?����=����>�M�>'kǾ�.q�48������0����>�*�>%O�>\�>�A�?�?�K�?'��>�_S?q�e?{6�>�=�'#?k�4?I��?��%?2|9��d�>��^-?�޾>m-���^�fAþʦ�?հ�^~�Q�q?^�
����Ԏ�Zw�>BJ����ľ
���*&0����>��?Y�/>��(@f��c�>�H�=g��yϾ�r0=��!�M3�k�~?Џ�=�>]�>]ڍ>u	u?�c6�[ip�u���܄>�%�>�@,�d��h	M�UI#?�*�>5A��;pD�<��?Y׵=v�о����j�м�>ݗ���
���W����>�h?V2f?.�?0p?�Bz���}����ܾ]�4��� ?w|��2j�>x���9V?�u�|v��W��1�>mGu�>�f��=lZ>��`�h�?R#�=��p�E��>�r��; �1�L?�-=��>1o���+f?�%�=O�տ�㩿�e�>�1?�-�e�:�<�?�2?B)�n���u�8�	h�?0ר���������G�?��[>�_�?�[\���@=�����5�i?3�>�@,?��0��'>�0�>��?>�"�N����%�
�!���$?�]0?j~�>�V(�Z�پ+A�� � �U�(�$X/��F��s�>DA����M�i��0>$I���q?*�B?�5�˓t?��k�2��=�� �%�<�5�<��><R,>�)]>�O�1\��1S�r��=��	���S���'>V�����=f?0��=&F@>{��=�y+>,�;�N���?C�>�;y�f�-�7?����5r�:�|?�ø>a"Q>P^�>e$?��M>?���M��v�>|>T��o=���>L�>.�>��*�����ki*?ꂕ?3�$=+�ھ�o�>�?rFV=����T��z6���"���m�I_��+���I"=")/>Yޏ=q���Wl?-H?[V�V��>��q>\��s<�H�=)?��?#�e�_��<�&>u% ?X��Ŋ���]��=‽Ƚ�w6�>9�^��{��f&>�ˀ?ϟX?B:9?n��>N�=���><�~<c ?�x� on>"Yg�9S>u����F�cd�<�?��(?�
�>�?�D?!O ����\ؽ��>M'>�)z�Y@>̰>�w4�0���U/=Z� ��S	�i�=;��=�>]?�uҾ�SU�љ��� �=�P?j�>ə���>��XD?�B>��=�k��j�?Q=;89�=�μQ0���;;���?�{">Hɘ=��ս��f?��>�ɂ>�\�>Κ>"�	>2��5n�D&?��?3*)?x@?�:?�v4=$W��@F?RN��V>�12>��<��2?Δ�>�s=C��>`w?��?��K�����^��؃?�j&>5D#���?a�?�Qھg�<��F`�?�<�=;��?!�̿���ˏf=��+=�g>M�=fG{=Qm�p*=�)��x�^=�Ge�Mvt=v=y�.=~�i���;e�>b��=S/�=�*d�X݊=a{�<�ӫ=�9���S�=E`=�p�<�ĉ�Bj�j���w�Kbk��}W;�O����;�d;�=�\=o����2�i=A睽�ͮ����'\<B�i>Po�=��e=�\>��%�:%��ʚj�@�e�j�k�6h =u��Y��M@=�~����;��lD�7��bd���d��f��"�N�<Ҏh��a
���d�Q>m�b���=����FC>�5>�7�=pU��`�=z�k=D��=�8�=xx����=H�=��=b�SvT����=�+��2���*�כ>�!>�.=Xn�=��=ec���6Z=A�R��O^�8V����6=I��-�߽������w#ʼ�>l�=\�>r�%>�A���e�`�Z�kV >k8D�~N���̽J�<Onʽֲ��)�������c�R�0L�
.���ν��<#!>�w>��=5�ȼ�����r�����<qyZ�ܑ���T)�lgC:��5=���ϰ��W<\�E�I�>E�=X�.>!<���=������&=�]�<��=���P��=�\P=�p\=Z��=��={៽z�u�o�ѽ��B���G;j�?:0uk�������h=��P�P�i�d�4V:s�ֽuC�;ĭ��Zx�P�)�Lק��<�{�)=�����{<&kV���=iV=�]=�[\�47 >)����>���ֽ߯(���^%���������=�m=�����@=�)�8���=-q�l}���\��ܞ��bؽ��9����CԽ����[�<0�Q=�%7=L����?�Oz�=�0�<<�R���]��%>�5'�d�[����=���<��,>с�=�4#>0�˽*Q�"����=)�c? ���2�dq>�;�V�Z�/���?u=�(	>�ּ=T;�>�#�=U�=��G�o:>{<jeν���<��p>d��=Q>�8�=w6�>%�>)ϻ1�=��5>K*E���=����V)>ɴ��j��c�A� �=��A==��w���b	>�N���=p��=�~�=�ݽq�>�i>�k!>�]��FF1>��=�Kl=�i�BJM�dn�O�-�.9.�3��|��KGJ�4�g=�Ѽ�u�����60�;��>,��=M�5���>z�*=�4�=~��=�>���=ľ�=L`�=[ּ�u������h��^$��)��4�R�9���]�+~� @3�&�i�K��=�G�=�2�=Qur� 9x=5��=�|�=W����=l&�=��;r�<�D�����ǽ�(���G��̻���<�A2>����\�U��jP>���Ύ��@���3�>�>��z=q��=��>��ؼ�X>���=�L>����a�w���*P>�@)��{n���=��Q=^�c�v�_�|*�:�\��F�=�ph��'=!�=>��=&z���ȽH�='�E��S�Z�Rq=�z�=*�V>$z=�8/>��M��"E=nd��N��=��>M��=o����;>p늽z�F��!�;�{�=��J>�L>�c�>N-�>�%N��u�=�&�<���=I�=����o_�=*�w���;�N<n��<M��=���=lX>��a>�gQ<�?��!9���='�e=����+�����=Mϕ��+���Sֽg��<O؃>2R>� �=��>�!�<�z >���=�yQ=�A�=�֑�how�^j�^�=blP=z�=�����PR�i3��D��g��h�~��tC���K�_��X_:��j���4�k����r���j�=�L�ד�=���$�S���5���<�R}=�> ��=i
׼�^7�-��=���L�>V�r<�>эi=t� �t\׽�-�c�����(�7����sZ���̽j](��"��r=ݮԽ`
�=\R��-�r<�sý�z�b���t�a恾5�?>�ý��9I˦=s�s=�u�V�U��'����=�!�B�{B�=o!X>�d�=��=g�>�κ=Q𡽧Ž|W<z�c<�#�֌���ý���=�O �[�����T���9>�r@>�^�=�>��U���������M<��=�T����K<f	�=��b=��-�l���Ϩ�=x��=L>�l�=�> f�=��=�3�=��2=֤=��"���F=q/<�w�=���<�`�=R�<*0��LV��M����=�����Y0��t��U�����삼��I<c߹=�\�;MQ�=�V½ض<���<>�Žj�z�R��Y׎��3��|�ȽK޽#�1�ĥ<Γ=c?(�B�A�� 9�!�<��;>�&G>=�?>u��=������K��䀾Cf�v���ν3���ee����C@�� �=��~��@=�BE<��ս��}�=���=+z�=��m>]@%�/Zt=;,3��U�=$�<W�����<==>�>�����E=:�>r���`�= D�=��<~���� =m��=:H>� �7>V��=�P��ؗ��)b��&ݽAg*�0�^=%��;�q>�/>�>��ɹ���= �m=a�=�]=�m+>S^�=�����]#��޼���K7{����;����Y�=��>|���j,�:�=��s=��="m�2�7�Ͻ�n߼��%��i>��G>�,>�>>��B>�qW>��Y>P{�=�<>W�>؜a>'�>q	I>y�T>y�V>�E>N� ���=���=1Y$>��n��^�=��!>oU�=�`̽�']>;6>�c>�<8�=��5���ry�@��aE���;�G�� *��:�0=��*=�������<[ӿ=�ћ=�ǽ�� �G�&���v�P`/�ϫ�=s�5�3=컅�qqi=�!۽ɯ�<�l�=�vֺ��=��l�=��o;Yp��Ȅ<����<=�=��]���'�����
�]ǿ=��:Td��u��)�!��໫Q;�'6��L>md
>�S�=�8J=j���ep����#�.��J�p=�=�=Z}���轢L?<�S�=�u�=�Խ�5��Z��e����!��& �h ��;q��G��=:*�=এ=�l����%�n�>��=�&7��@4���:I=�<�����~�8;�����<w���R�=��=�~^>��a��}J>��=�C�= Nt���=Yr5=e��<���nV=H��=�=>r�ý�=�:�<o�����F���j=6�ٽ��=���=���=Zn�=g?�<�Z{�V�>�W�=`�J>7y$�Td4=ɠ�=ǋ�=�5�߄f>��>۹�=J7_��kV�n5��۲��
�  >t�=/*>w�:�>��=�z�<�̳<�����Y>;o	>���<�(�{֒�D��dC����s�(���H�:i"<���=��==�U�S��=�%���躩(�=TY=�b>�"Q>P�L>+�q>�
�;
�K�ؼ�1��=)��=��=�so�\�>(�=W�;���=,��=Ḱ>UF>�t>���>nb�=6��=+L=����_4�=���=����H�ͽ�r(>9��=���=b�ǽ>�����P���0�Īf��xɼ����'/�>�6��Z)�B��<���=���;��t<��=�{�=Q��3$��%���
>BO����(�Q=�2E��s��I�=�$�=R���%=�HB��9��:ƽ4�-����=��>xM>��+>�e>Q�=��2>Eb�<^�>w6нd ���G���<=���u��wJ4�0�:>ڑ�ro�A�4�<�9̽���<J���UGN�y�=�)�����i�Ž)���z%�bbX�M���Cu������;�ݼ��ż�p�*�ؼ�j0��c�=d��=�P�wԼ��U;��+>$�e�w����y&����<�н�
T��*<� �����*j�ԫ::�b=������P�>�d�=~�	>?Vw��[�=��<~�=��>��=v2>��>n"|>�="�	7=�"�祳=����M����%>�.�;]Z,��S��I=��-�@7��km�A��={Y�����M�W�W�3���:��O�T"�K�=)Ce=��<n5@�5A���?+��o��>�f�=sh7?�Z�h��>!q��&����>���>��u����?�_o=�B����>�RO?���?�K.?�+I?�����5���3M�݀��\��%�
?��#>��?�t�ʾ��n�B���Ϯ>����7�[���G?П\�S¡�=���"6<?P�>�㓿~�s��z?g�?�^�>Ȃn?DP?@�9����?tǱ=iԛ>�U?�w
�V����>1憾9s�vk����l>H?2%��Ǫ�>���>|�ҿ8G�)����Yܿ�%��!ג>��>�I?8�ۿ0�>�4?h�f?	���.@�:Q=Kx?�d@?��)?�7u>���>:��>\5�j�_�oY��>��>-����`��;򾄪�>��>1�^���=�y���׾S����m�����u�L�&�=?C\�?ɵ�?����g��k�3?��?W��?���?[��?3��2Ҿ��3��9�>C���]��o����H>+w������shG�t=?�����7��gz¾C�D���?���>��#?-a%?���=|��J(߾�M׽Fc�C�����˿>8]���z�>iX>³M�e�i�P(�?�Į��x�O����s?���#�?�^a��l̾�ش>�,=̬�$�R?X�@?@��))1��Y�>*��#)|><+7�>?'9)?���=���?D`�>� �����>Mt	�P¢��Um>�Ys��Y���Eg����J���}1?	��>;[�R�C�>�>N��*7??�K�=�1@�{������F�&�W?hI?� ?TIÿ;&{?]?��>^�f��;(��V?�x{?�%�s�"�\�?����EP��d �wBR�o��>m'y��<�����=	\Y?y����yB?�%7>A�>�:Ѿt�>�4�?�X.���yA�>�X]?H�?��>�d�>�*L�jB?%���<�>ll*��Ñ?����f=?��+�
=���l�B=�����7��/��?.*���P���J>�7�?a�����>?�x?N�v>�혿��>��?�F�>�;"?��0;	��ꔾ>�k���:\?z�*==M�3%}�y_m?�c��;J<��>��L>�����?y$�?s]�>��A>���?��_?�!�*�?�e�>��?�ο0���iH�T͂�	r���ǔ����oʟ���ο���<0���!�=�S����?nd�>�z?�^ܽ��n?WQ?��X���>�^?F�Q?��=V�>h\�XǪ�Ïw���<m	�>_X�?a�)�y<� }���{��P? ��>���>x�9����?>F�>��	?V��O�T>�M?t�=y��?�i�L�>�R�j�*�g	>q?6���V���-?]�d�5���\��O2�>� ��m�i�CAe��#?[>�sm�����.�>_.?j�#?GH?�/j>ː�>��^n��{g��h���۾4���250>@s��Y���0��<ھ������o��=QN�>��.����=,"�T�6>,t�>$�¾�u�\��c�;>��ɾ7B�>7�>ɶϾD4?�(��Ц�>:��!��e�>�e�I��NBG>�� >����:>�=�>q{ѽkO�X)�,> ���:>���9?�ec?☴>Ҏ־�s>�}���<��/��Ѓ�;.�}�/����.?�!h?q2�>��:?�D�w{>���t����x?ҩ(�ۍ!�N���,)?���>�F?��M?!v?H�>���>��>?�-�H���7d8�� >>1��>�>H�2>�ڜ���L�����T����nP>0!��>VY0�� >%�W�c�?��?�-���OS?���1@q承W2��L�>!�'>�i�&��>*v"��d@@�?!�<�
Ѿ&�H�I�о�:>Yqc��t�QIͿz�����?�־�-<�ظ�>�̉=6�K�J;Y?8t��ǎ��}W> �>|���I�>�	5�f��,S�=l6��DM?�rs=��=>f��s,�>1����`�;�  ?�$��pf���H��e?�z�=�������>��?֒ӽ��<)m�����=-֢��K���?���t?:ʻ�~����~����4?	���ٜ��e-���r>�XE�l�.�w"'=�H ��>
��;�>�1(?r��������o=�r^>JYн/��J�ǽ�Ǘ�����F@?��?�gq?ڟb?Xt�=��*�|*��|���ʕ?�>������f���Y�ĿiG;>��ľ�a?½-?�|�?e�����?@��@4s�>��#��M�=cU	>��A?�8��[kf?F�)>�.���jR�$}�����D��W�J�|	 >Rg2?M��>���̱�?}~?�FƽT�'=��>&�\>�����N��j >��?�+>����~�=��\�%p���V!�s�?4K5>~!�E�]��>�@X�p��F��?�ʜ��N��%��=���?nE�W����r�>[�?�=M�-Ʒ>Nʷ?�9�ҫ�>z�'�'�?J'��(�?&3����>	�"�uݻ>�Gs��W?]�����>�E������!?
(B>�{?�L��@X��?L?�>&<?v�kK�I�����>�{}�V@�x����
Ŀ��>,�>3��>��x� ͔?a4�>*�r?鐣�D$��?��b?��� ��3��=�N����bl-=�?����:���۽uy�>�a?�O�?��<KQ?u�,?�v	>{B��ֈ�??�մ>�>pδ���>�e}���P?���0S�?���>�><?��m��3?����>�=�~;�Ȳ������>���U���=c<'�����=h�>?�I=��}�[&?��2?:cD��8t��ܓ>��><���xq&?��>q�>�;��?���n>n?�G���R@�f�;׏���=C�p�ۦ>"�X?��S�ֶ�8ս�����=�7����E��:%�M.?K�^��E)�G��H�?��G?
h?�Q�?���@�?�T�=��W��z�>���?2�?�����2�>�˥>�3����<�s����>�t�X�)��G_?3F�?��=�zDǽ@�@�8������}��;2�?�{?'c>���Z5�C���s2���Zƿ=���aSo<�K��ʭ��]�>�>���>C/+����?��Y>��?��ſ|������� >��J��B�>H�r����>fn?��o�>������>4ӊ�[Aa� ?=t?򌣽�k�?�[�< ;���� >&��l�Xe�?5�=�[�>�Q?�v�Ay��\ξ�����>`_��&>���>�&}��#�= ]�>�%�";\?13R>�?�?�<?�ܙ�Vk>$��?�\3�6Չ�� ;�p�?�*;�a��BC�>]Y�P?�9�>�Gl?�ZV�q�?�'=?_�7��+>y_�e�0��=Ck|??��?�3+>e���:y�n���c��=�/���[>��?��?W��&�_�)��BI?��S?B�?Q�D�d��j>i�>Q��={����t�?��>��>2���07W?�R?��>B�Q��a��������I
��R��}�>��>����3>=�?��ɽ�}J����=w�?�<�?NvK?�U�>�z�>�+�>�X�=�GI��\ � >b�G�H>�vڿ�xp���1�mܙ��C?�ʣ=ox[���སo?��U?K��>R�@?��?�G?f�>�3?�1����>� �=`g����?�K�=ES\?�jx������#��0[=�����2>
nS?�Q��騾�u>�"e��������YDɽŞ�?����;׾lq�Jc���;��Z�Ȭ>M��Ռ?�0���W?^{�>ڂ?b͝>��f=!(T?�h6?�3�>@�S?^��>\�{&?Qg�Xs�W�Q�S���H�� ���uƻ۷>�4��Ƽ�>/z�>�(��OtD�P*W?x�>ϼg*?@m�>o�?=]��=�w�;�=��\w}?�Ǘ��ֲ<0�?��?6BT�V�4�����Z�4��=t�>| t���@��A�@��=0��U���,M�eNz?�bm������j�I]@�_#>��>?��>i>4D��ev�=�YD��N�!�;A���Fm���>�N??�r����?���?GA�7��?zi?�\%���^�ŭ�?�w�=�8>�e=��?hv�>�?��5>�s����	��!�>���5$��]ߠ>�&>z���]�M��?R�Qˣ��z>	�h>"@f���>������7?�\#?�":�\~�$ ?(�D��R�?n��
,=���>�c��Ń�Ҍ?S?׼�Oj���>�i�=�!C?�n&>&uP���&>��о��A?���s�=iZ���>�k�(ML>��?&_L���`>�)�<z�C����>�u�?(�?6ec?�ӟ? z?e@??�.ɾ6��<�#�>��<��D����=C�>����n�?�MƾT�վ��>RV��mt>���̊���������z=�L��?Fg?_�پuQ�>�V>^S�>�P��!{O�r��=�放z;����"qY?�<�>nK6��,?7�鿪��>%.4>Pq��*�?�����8�KX?��|�vۂ��=I��B¾l�B��?5�u?O�B���A>�A0>�jݾ, �y8$��`?�?{�?^񒿆�? o���7駽jx������d���+��?O�'?�U~?k�> ?0Q�>?
����y?�T?d�ɾh瘾��'���\<�*�=�&L>��>��¿]���5��J7����>IiQ?]�̿���?f%?^������&@���^��,�>��J?�A����x?�L>�☽?E?���>�6�>b�Ծ�5�>��p���q=T�?n�|���F��5�'"�?����?�#���k����Uƾ�L?�{�]�c?E��>�?|	@B/V?�2k?��_�c�=?�nտ��#?��tU�= ;�>�֦�R�>@n����ֽ$���:@�<�ڼK�>l��p�'?��d?7���|������\�=��!? d����n��?Š�>��2Z�?�� ���k���q?� ������[�O�;?e���?�@�=���?�78��&z?ҥ>>�T�?0H>��Q��A�����-�>�I��3?eoR���?V9������b��d�>m���R��?�9K���Q�
��������>���=��?�;�>r���P����y��i��>��!�2w?\�O��?����w�����?%]*����&���������!cɾ���>Y�=>C2��6��=r~J�>�s��C�=X]��^U?�=����?ܘ��Jj�?�K���Y-������[?6�|�������1/�>z������-���,?3�P�d�J�1~?�"�?<�>�x��&�C���?���
��>�����($<f��?�1�?�<?��?0+�����Ψ?W"�>��;ƍ�Qk�?�$��>ݔ��#��]+�p�.�݆*��!�V9?��G?���?�5�?�X�>9(?P��VI>Z�)??Dǽ����z���$�U�M�'����D־��[?�Ͼw� �k?�)���S?�c�=�˖?����\ @~Y=�¾]K�A�>MP����?Ί���9��^�0U��1>3���?��&��-=�Hd�^�U�:�$>�F�����z=�W?D k?8�>���?X�?�	��ִ��H���~?���x��<f.��<?C~��9�
@����fK�>a���JV�Gh=>}�2=�O�p������[ݾ��<�J$����>3?] �=���>����b�[�����?�(@�/>��y�������?S��Q�>����ǌ?9Ia>|kD?>���w���`����۾�!��d6��l�>X)?q��?�*�>#R�lH?��˼x�I?t��=j|�>�Z���$��W$?� @��>Z�&����>�G?l�[?i�?>~�>cEP<���ʑ
?�/���h��� ��$> }y>���a�'>z�,���>д�>J{?7�>�+w?Ů�>?m?!岿!˿���?�2��Ƞ�TX�>p��>!G�>�Ĝ?6֚?/�t=�u@��'S>�N\?ue �{
�UX���V����]�c?�׽�O0>��説>��>I3??��>�����J3����ë.�#?��Y�Rm7�Z�2?$m�@7���f?i"">Ѯk? ���c��>�/6?��*?Pp�|�������?�?�ܲ��=�>+7b�.����'���p> ��z�=��,���?���K�=d���[?i�>���>u'�?�\�?��>�d?($�?5�M>�*���e�=���?ɴ�&/t��ϵ���>���=�;�>�o'?���� ��?t(̾���_H?iF׾���>i��>`�Ѿ�_A�!�W?�dG�r��N��>_�@#�>cќ���Ž��#=R$�<�7�?s��?��=>��<慾����;�����>��֡�;[����v?Ȓ�f%p��^���߾B��� ����%?<�L��hF�9Fg>���>ӆ�=�.����<�� =��>3c&�!���+	��v��O�2�j1>>L�:?���>�g��SM{?Q$I�L�*?�::?���@�ſ�>�m���?�W߿���>o�>\��$��=��k��)�='��/j�>�3�?���>p�M�T��R��?�J�>��>A�?ݿ>ʱ�%oU�����\?� >p%h����(<�!1?��12�#h=>�?w�E�4C�x�m��!q?��?����������	=G7վ>):>�f#��s�>�U��-b>�U�^�7>ek�<�L��D?��*t<8o��dcX?�X=�c�>cԂ��^�>f��>Y�'?c�ҿ���N?d^I?�x��.|?"�?M�M���P����E=?t�?`�>�)?"s?.i�?��Q?�?�S�>�s?*�<?�� ?�X�=�0z��w/?>־�쒾(�?��?v^�����'�W�|�/�?�݄?��ľ6!��hؿ�8/>��]=���[c��i>��獾K.>��>dy?�X?��k����@� �>lI�Z���>�$���=�=�>�i�Z���)G�>&~�>����|�?��?i����=g���>��'?\Q�=���3;�V��}������Ayw?���=�>\@?� O����>�o�?큤�e��?�-?�=/���o?����1�P�n���?�'�>0�>������B?�'���@���M����p?'ʏ>68@�\������?���>��?ޕ��]?.bſ38?
4"�������>���>`A?o��>��>�x=>q�� ?�����Ӿʬ�>�>H��VcǿiG�=v�4?�� =�> %����?Ź(�_?EG���ɯ?ͨ$�����\
���u�"��>롓�2(>Gb�>q�O��<�3��j�>~�?�vQ?ǐf�	�?�᡿�}���j?q�&?���g�i>[��$�Ծ�?)�?4��J��>?�e;�1���r�6H7?)�ο�?c$=>d�l?��7>h/�=�R�;�\�����>\�-�O�?���G�;���>�g?�jx������X��o>4I@�e�?E�C���?c�ÿ�S�>��&�k���8�u�
?}�>K�@>3	?CeH��`�VS�<��¾�d�gYu?�&�憏?���XZ2��̌?cqO��β=��.�4R|���n?x��>X��>d��>�x@?�⾤�п)2>S��>L����;�ET������*�ͅ辺�;�>�X=�E����c?�14?����4�*�`�n�V�~���Ľ�y<>*��?�N�>N��>k�<uT6?�Iݿ읭�v�+��N�>̪����?�� >}#�>��������n�?�^�?U���]e>vL"?�l`�m ^>O.>rӨ>\�N���f��Q��8?��>��¾=�@rf�Fn�?��>�Ͽ��� >ދ�>���p(��]4?V�@���>��Y?n��i�����W�j��=�A���г=ꉼ<�wþ��>��F�ڮ�w��?68�xg5?C>��$��?�<8#=���>x�C>7��?�HL���i?l�A>�66?���ҥa?�g���,�>A�>��?�/����*�>#�@�ф?������ e�R�>��>���>.4׽H᳾� _>�u����<�55�k�=x 2>�=�>U�Q��h5?tҾ$Vi�S)�=
�=��>t.{>�4>*��>b.�=�r?G�>�j�=�3`>2N��lC�M�#�ˇd�n�=s���><�ݺ>yU�!�ھ��������ni�Ī*�Ly.=���>9>�n7��?e�>�kF>�.K��jj>I���d2=W����#��ӛ�:ʱ��%�!��>�VC�헂>q�;�X�>��~<�eQ�Ӑ�� ����U����"���>Y�=�O�>C=��Y���%�=��>E� �is?���=�i�>ȵ�>��۽�W->���>0�C>��g�m\���U�<�<����oU��>?c��/��;���Q�>���>�xW>x�����<�t)�����/UO<�S��uf��/��(��Ъ�>��?J\�>��?l�?��p��H����>[ =p�f�&u�=��%��<�wI��.�n�_�譑=k]=9=?�ؾ֬��<?�>� ?�?}8�>��>��Ͼ�����@��v�>��=8+6����>�Z�:�d&�F幾���޴s��޾>��>jO�=��<�Ծ�ͼB�N��Ř����U� �O��>Y�?ݞ�>�~?:�����ӽ����jؑ�D��/��=���=G��>�3��*3?F�!?�C>����b���<�\�����1��>7x�>^�=wD>z�ٸ��՜=9�?>Du>>g@>#�n=�(>�>h;]�8y ��Q2�T�>�����n��Z�~��<��޾߂=d>�?�>�>`]>�֫�F�>��6�9��>_�>wT?�0�>M6n�^h�.��e�&�Z �=���>��>*p>�? -?�t�>o݌��u>��>G�>���>�ه>�>�V��io4���>�$��_��=62ƾ��>�9����w��i��c�f>d6<��= �>.�=���s����?��K>0Ӆ�8��RE�>�	�PH����>�\j?�&��p޷�������=;�>~�>��R>�����I��B�>Z����=�o׼j�=׿?�j�j��F�d�h�>\�p�ng߽�;���>��o>�a���=8�)<�A�>q�پ�	=r&¾pA�>e%��ϼ{%<�����Լ>����5����=L���>�ϼ9���t9>F~Ͼ�p��Y�y!�>ǌ�>��8=��>�+\����>�ͣ=C�G=�Ě�d�;?�D3�3����" ��6>N�b��`þ�G���Ė��H>l��>�O������N# >��G=�@_?����_־�8�;g?�1�=�K���T�&�_�A��= �
�d������>+B>k���`�r��=�rݼ�F�����W��>���B���$>�f�>��s>ⷘ>���>�W�>ʈ��h�0�r����Wx=q|Z>���<�N�N�>��\�^ϾC�C�h@���u>�i�>���=򻺽�(��R�=_C���r�9���a>��J=��<pO�>�3Q?�\��m80>Xٲ�ȚϾ%d��6�9�>���>7�>�k%?���>,�M=��>r=���ҿ>y�S>��}��6q���U�쾵��=�-��Z�^=����bw��`?�]>VZ�>X�?N����T��(�����q>��>�[>0f��8��;խA=�_=�(m��
���B9������w��ξ����K�!?>9�>U�*?T3k>���=\���L۽�s���8����>'��>�ڽ���J��=hz���ǣ�����A^���\���J���ȽB<�}ހ�!0��á�M���"��d>�"�s��щ�i�>w�� v� ���6�`�&󗽖<�=x�v=���=E�=^Ö>ð2>���<Ϻ�>��>��f�������ĥ��AI��wc��������=�0>3ü�=�y�}k뾷-|>P�?�Ò=��>�_'��`T���徊��s0�>�)�������_<�I >�E���m�'��x`�܈��P&���콝�#>��K������>V�>;(���D�`��/�D=��+�C�߾(����<=��N���	��ા��K>gd&���=d��=�(>�#ϾSA����>yo��O��>��?D�=V���#i%?�祾�>#�>��ɽ@��>���>�U�}.>��5>�r%=^�{>�N
?g9�>�-�=~N>ǳ��쌙���ܽ��7�������ʽ�J"���>�->�I�{�p�8��>���;<��>kX�>��m>Q>uT�>r�?����]�=Gjk>�� =�z>��>���>�S$=ľ!��>��<�^���gL>�U?D�>圕?���>���T(˾T�=%~ɾ�(H���ؽa���ߺ���S=aH ��}.�8L5�S9���.=z/,�s�����m���ּ�^>�Vf>	�=�$!���ӻyM�=Ā�>��S���r��:���;�6�/�s>Yc�>�O�����A�cb�=����9;%97�p�>V&�>�����>�H?�7�V!���C꾸�8�C�=-��=�>>�S�=��*��k��x.����=)���(ѐ=�dQ>C�D={���yͽ��w�E8���S����aLm�h6�#i=kks>0�L>Yr���ھ>�??��;> g
���>��>̏���l�d��>q4�><d�>V�m> � ?;e!?�^�>�'o>�?'�?�
�>��x>A�?��"?��*?m�r>.h��%�%��d>L��=���ݥ�#�{=0��>���ɮ�='?�=qH
?s���3�����=��>�r��'5<<&��+6쾒e�|"V>��>��½�=%	�>��>����,��'>�3署�Ͼ�">� �(}�<ώI;F��>�i?Y�����>ܰC�P��>ᓄ=�"����Q7ž�&E��b�>� ���r�R�(>�e>�N��
=��Ǿ�!])>)�&>`*Y=��`��i�!�>3o/>sĆ>l�>^>�=�m��a=�����1�˾.���qd��=���36_�G|#����iJ��yw>�ȍ=��47Ǿ©l�CQv=:�=>Z�?����=�E�>���=��>=��>c>�>���>M��B�=ll�>��D=㷒����YR��+V���>���#�1;��>�j?Ul��W����>��q?�s�"�>喼>�?X%7>HG�>x[?b&�>7��>-+ھ�\�>����}U�=�Ѽ�ӻ>[!�>�^�>���m1Q?R9��;5��:e�=�d�=c��>�R�6�D>�P>��?T�y���=�&�>��l?4*Y��D�=k����>	kM�ߺ���<�e���h�8;���?�>:.��v���!%ž��>Y��rl
���;�[оL���Y�;:���,�=��>�,D=�x\>�ԋ>P[��j;���8�>�E�,�>�q�;���>�`�>�)��r7d��y=XԀ��AO�6
�=�W(>��P>�k�=�ƾ
���t�5=��>�?ـq>���)x�:�<vk#�/�� ��>�8L?��^��<�8?�\ ����a���qY$�?��}@��Pm��C�7#��~ɽ*�> ?�?	�>z�*<d-�>}��>颕>���>8ߟ>�z?��=a=}7+��b���X�AV�=�>й�>�NU?��
?dC�>��>�>�Ό>7԰=���>��B�wf�>63?t ?B�?�>Y����p<^5����>�L���R�8����^�>�L+�ĝ�=�u�=�y��,h�v
�xz���f�m :��݆��& �>婽�9�>D�l������(v3����IQL�p�;?Ѳ�C����62>������=P�;>�@�=���D ��N�xw�>BK��6
�@㙽��p��.��� m�c<^������ǾK����H>�"
>�%¾�&_�_{Q�q)7>#����$�>,�>=}y��81c>�=8?�g-?��?O!�=�w����&�>���>�f-���=IP�>�">b�}����>-B=]�?�V�=�/�a=C����>��b>�0�{U����?��辰П�SD�?��齬־�����B��[d�kD��ӄ�9�P��h�1]����LR?x�?�~>ı�=�M𾸹�?��D��\��@*��*�d�=�����ɾ<��ZB�>�4?��_?�^S?w�?ǫ>���?���<�ŀ>Rf��Z�����RR����f=��1?)>3*|?qa>�ϣ�r�>f��,4���־>m0��0_>Ao6?#E�?Ee�4�ӿ���^w��(�T�ϔ˾�O�?M_>aF�"E\?xh�>�\�=%??�%?H��>�Ԕ��}��$q�jֿ��ƭ>�1T<"^>�����L?`푿�b�?���?���?Qd�6 �a�6?��@�eо�?	�LS��-�>� N�U+��C���+G?��˾!#�k�s<9T?�M�>:��>���?V�N�T=����>m�>�:�?:� ?7މ������l�{����*��f�>��E>�/W?t�@hs�?�0S�/���p��l��@X �?�=�<����?/�=y>�?J-�����1��s��?�q���$=�Ӿ�%X?�����u���r[�ʆϾ��>o?�L׾�Kz�we�����tt�>~��ynk���>:@�	����2����??\b?m��m���PO��Ϳ͟�?��>L��5����CϿQിjv��&�2?��>!֥���>�o�=ND���a;��J>%�?�(9>C4�?��|? �b������>1�?�z�����<���>9
��L�8?-)?�:?W�Y�e��>��'�x��>�S)��&��.��>�s��:�Ҿ�n�>Ż���!����?䄻>��>Χ�?��?Db9�F��C?
豾�
w��7�?�h�>Ś?��5>�{>�*��G?�������^��R�3?=��%��?7�Ⱦw8�=u�H���>�<�>q��?#{^?�4>$��� v��0!����?�X�����=k��T?�?�M=�-z>��I��� .���P?��7����W�V=Nj�?�ޡ>!����?��6?��?Ŗ��	�<ld�?�>��zI�>���>ٹ���½t7ؿn� >��羙np<�vn�rh��C�?�.�%�?�R۾ R�>�&�?�&?Xg���:?�H >%��r?��>���>`���e��?�-�?�%��%Y׿6�A>�S;=q.�9=����7���Z?1�4>�i�>���?�4@Xc>7�?L%`?Ŧ�>+@��֙����>P�?!�U?Д!>c��><E��e3b�-<�?�?㇩�}p�݂i��w7?_翛��>0R�?�-����Ŀu�\�z���Q�>��>���׽�'���?>��?&9�>W#?�?h�޿�ĺ�<�����-?l��>錄���>3�+��M?:L���3���>���>~�>����^?����I�l?��Sv�=V|>O��?��?��5?���?_^o��o��5�h�sB׿����Gu���9���Lk�xwu?D3A�E���N�>W�"=�p;>0d�{�.��?�>����"Ï���>O����V�`l��z]�>Q�?ڠ��7��<���=��`>�ڔ>K6>�L�?R?�5��?���׳���E=^H�Pۺ�&��_ 1>�?h�?{����"?z������'?�?ǿ�>>��?�R�>n�'?�y������r��V@?֤�?���?4��?�Ŀ�٨��BZ�䎏?a��<sY�=��>��?�����1��.[Y�Qc?IO�>�YN?}� ?�2
����Y ���hu��)�=��=l�=S����1�>�����b�R��%�E>�W�?�y����S��:R=�����2�;NZ>����9�N�P��>�����p�iM�=b���P��?H}���;q?�����@�>�?c��?��?����� ��L�O� ��C����x��?�'�?�8u��h��P�q�n���^˿�>R������>���Շ?�,>���?-�?G�:?��"@o�?����>��:���R=�'���ʙ��[���i><��O,�.*?��/?Փ���Ŋ�K#����y?w�?���>��&?�q�)���{Ǿ��a���> �>b���L�Ǿ���>H�<���˿���!�?�\?c#�>|�>�s>��]����X�?�
��ƪ`���X>�g��5��b��XƊ�~�!?m�%�����{?ȉ�?}7�?��?(�>4Z?�����?�)~�����>�Q�<�8�>듬���ս\��A%`�{����5ʾ�,n?��B?&n-?0��>�!c�X�?�~��rf����>�H�?����^>0���rC|?ye�>,[Ŀ�ྶY7�?� >?3��?��?��<ehD���u=���$2r?���?���>��Q?��K??��?��>�(��o�/�]F���D�e5+���=:|�����H��?R_+?��K?���>ُ����O�������?�y?�}�14Ҿ٭?�V�?�75���3����=�2�?�S?C�� ʾq�?9,'?b��=��p6N?@�@��v����?\xv�z >�&���
O=sY�?ݗ�?D�]�_x����ʼO �?�P���n�>|*�?�KϿ��9��y6����^?��?��	@&Nf@k�o�=ͣ�(<5�������>2�?�!�AJȿ <?W��=�0�>&\�>EA�>kSW?�۬?W�F��s�?Ę�2�̽)Ö��B?�i�?A��?Dh�>=yX?d��?	u @v@��M?r>׮�?��>��>�%v>j�>v���Dg���?e#?���?V���H�� �>�V�?��
�ϡ߾6�,�0�?������q{�C*��L���+�>j?n�Ҿ�L�>A��>!r(?@*��~�v�� ?��>��ýߜ1��:�;�*�#:��t�?NP��%p�)u ��~X�=C�3�¿���@/�vR&?��=�O�q���.,���Ͻ�/@V�zjH>���������?tS˽� �^�`?	�Z=.Q.�����տ�>�\�?�?Ʉ�?��?�>úM��7��X?f[��<�Boq?f��6�?kM=������;<��ľ�G����5F�><�m=#a��Rk�>
��>"H�e�ξb.��Ű>��?�V�>�#�c�B��k��|�[=�O�=x���l��f�?59�?~�����?kA>��>��rP�����>>fK���=�����?����<�?�H�<�?�U?Ѓ��=��i?)�j?�z�����4t�=p��>�䧾��i�M�����.�b�=�M�>��4��վBւ��>������;�c�>��{?�a�>�c�]�7�>��>;����=�=A>:F3�̲M��ID=���?'��P^�uV?�����	�V?^+L��A�*��U�&����?)֗?=Lk�q�6���^���r���A�;�B���q�����>%E�?��!>q���
.�?�Q��Ǳ�?��U?���K�gC��V<H��4%? ü���ټ'4`��>�>�BX?�#A>�X���?2��?]��?��5@�`�?R����� �>뾞�)�8��C���E?Q�>Z���Ӟ>R#�>V�(?ɰ�pj��TQ�]޾JOu�oC��i#/?�U�?/����t}>��Q>��=1�?���t�?��a?�_>��Z�?�[@n�?�M��?��9�1�ƻ���>���>@
?e����V��E��>�ƶ>�����@�?�?yr<<��=t����늾s����#��諾��>���a@n�?L2������.�7?#�F�'��md�>��?JGO?1�o�k1X��ם?5��p(4?6^*�2+k?C�?��r�E˫�j��|��>-V������q�s_�>�?��å�?5�mE����@��6���^?���=DІ�JQ<��y��~���k=#��>��q��H�>�?P��G)w=h'�I�G?ǣ��ҁ�q��) *?I�?��?e4I?'
?�?���?�t�����H�0�R�>��ڡ�{
����)?�~.?��[�ZO�?�Ѽ�H�쾂}g�� �qz�?Yӏ�v�r���rz�=� �>@��u�T��Ɗ?%�?�y(?wѿ6U!>8[E>o|�ʐ���x�L+�=��)��q���?�>ԭ$���>�ǫ�љ�>�oV��x���U� ���l��><-?#�>˟4> �=?���=�,�Z^>���=�=?�r�<ԱU����kA�4YɾBľ��?˿��R���|>�␿��\��4+�'��>������Q���
?őQ�{�>�4>��=_k9��ۤ?~�.���N� ;S��>�ľ
����R	��j?��)��'����2�!�&?M��QL1��%��S�s���Τ���E4��x�>zU%��>r?ҽ@f�{	>�F�>?�nm�>@�>�a������Í��0>m��b�>(J̽����?a�E�\��h= �B�A�e�+;����>B�%>R}���=3/x=w��>ܲ�w%�>�{�>At�6?T�d��4'?���>�B�%с=Y|�?I?%?;/?H�D?oh���4�������?��2��HX�����}a�xͰ��)���Y(�m=?�߿?)�ʦ�����?h�>]x)?�?!&L�-?� C�bۃ=�� >L�>?�`r�観?˝������e�<�">�L!��}?@���"]�F���/�>I�Q�b.?���T��UBr�|��>��>/O���4>AyѾ��>ܖe����>xɾ)��?c��׏\?������}���?��H�=��<�}=EM���@�=�L��b<��t�+D��>���@�>A��>���>i�>9�>�־�y����>�d��cR,���ʾ�ք?ܯ����=�&>>���>��>��%?5>�QU?1,=��H�~	���'a>��
�#�(=Y-���޾5(�/��/�G�Y�?�%�=L½�h7��>T��Фʾ�6��=?6�>���=eq�>��>N)>��4���>65<��о����9�e>y8>�z��$.�yl>k��>yMQ��	�> $k?ݲI����H��?B_�>)�>��U'>�?��>M?�t�Y}?�?��7=S�=�Q?v�@���>��.>as>�!? [�^���O�:��A�>�������>ʲ�=�1�������ͨ���-�,|s�f/<ۀ�=Y,�?й<��>���>�a���*���1�>�-s���o>@�E�S`�>ޒ���᝽ ���6;~�.hM�DFK��C�����.�?���n?J�C����'	�<�?Y�f���V>�=Q�h8���ɒ?�H{>���-�`>�x�>	�6m��X�>T�-�4�:>?Ī�П>�L>c����&�:����?�︾��?(w��I�>v�>�b#>�Q�<F����%����=�UN�]O&>g�E���Q�}��z� ��3��#�?�%�>�ڽ��־�[�<`�ڽ��M���K>R5�>Y�?4�⣪��U?��?�iR?��?�d�=+G'���~�āþ.P>���>�k�>��>O������<^�>���;pu>�@���t:?�x�>zޯ.���w3�>^����u�^�?��>:�ǽ�>ྉ�w<,�?�i��<5���>]>�<�=��4��#�>QV��?>��0�Z]���O&?2$S?��{?��z?RZ5�;���`t��^����?�l��G�>�m�>�Ϻ������4�Q$ͼ�4?:�*?y�E?�W?c��>
�T�]�>�X����<����;�=ƟC�W{-�;��B�=�y�>��
?�O3���?���>}��>��=�4��q8���]��>k��>��T?
��>���ؽ&B���ˑ���D>��>�w
�	�H=��">V�;��l~>NF?����0��&��kP?��x=���R��>�6���Ὄ�=��|=ܣ�����?񹟽K���r0>�C9���<X5��2�>�Y?<�`>��U����������{���>G�$��0�=o�=���w �?#��I3"���=<�>�8�>�l�=�1�������N�|�G��>�q���$�>���7>�ľGE����ԾM=kϯ������J[���3?|�>��'��P�<NU�>��>��b&���g*?<�,�������t��

?�|o�r�B���G�iy?:�>�HR�i�S>�_�=�J�\�h?Z��>�����v>��<�?�rc=i���0?���>�.f?���>��H?�V�>�l?�>�F:�>9">g��>U��?[a�<���=m?�X��2�?���>Q�b��h-��$4��J��jӾ��i?H�G?X%�>��(:P��b�*?|+�>l?���>�[�̈�[FR�u��\�>	�����Y>�?�l���Щ>��>^�`>��m>f��>>H �y�>d�>}hR�OJ?�#�>PFM>��Z? ��K�=�xC>ќ >?,<>N�Z�`��=|:ͻ@񇾊��=R�
��p����l?&ǽ��R�>3ܭ=�m�������¾�}/?	�k=�3�'���1�_>��<��L�7��[�H?�?"'G�L�=>���>ү�g@��A�>��?�c���r�?g�=��=���j=���>���=��m��FX�E��x�@8�>��.=2
K?L���س�#�q�I�y>��>:�>5����q;?.��*��4���=�����G?	m�?�G��*�ut�>v��=�_G?䬗��_�<F
!?�!��߾�r>��>��6�\=��<��>yC?Ge?x�?)�?���?ŝv?���=`�?��>O��=��/?�>��>Y'->�Y���^>��?��?�,�F}���r[?���>~�����8���>.�`�"�����<q̨>�����:ľ�f��iiJ�⣾�x[�bJ�>r��>u��=舾]`;>wmW>��u�<%����>�q����u�f9Q?��Ѿ�!f?�<?9��~l@�]kE?�B��X��>*m>��.� |?���6����T�>�T���X�0��=֐_���>��>ȏ��P�������~|��Sľ8���C���;?#?>ʆ�>dVr?��=��?�d�͈��N�m�dR��m�4?�ւ��[>�)>�w�<&�۾�m��~����sM��[ύ���D=��򽾔(��[޾�N�?�� /�=t����=��>	`�]
�=��h�?�Љ>�HZ��g���#?�kb?�;����X
?�Z�?5iD���L�-��>���]�wW<�/Ŏ>FW����>�F��G����>���_�>>�&��R�5:Ⱦ������>z&�>��;jm!?�#t�S3%?��̾�t�����q?���$�:��t�<X��k�� 0��>u��=3h`����-곾�>d���%���>JE4>�4�?Jv'�{��>�)�>�s9=����#S�<��Ͻ�ۘ?��m�
�+��U� P+�h�Q?��(��pv�D]e���>1�ͻ^d:?4Bq<��A=�˚<���=�l��>��V$�Y�=��=ut�>d�z>/e"�E8˾)���r]=��B?�O>}Ui�Wp`>�����?�K1?������>d�>cwk>D$�?�}�>�
���8�>�$��qy?\a�3)z?q�>� ?�=V>���>����t����w�0?[�"����I20>���>,ʓ>��?�恼m�L�/@V�&�پ����*�>L�5>f��ȻkbA>�#��^m?�y�����U�=;+ݾ���> "�=mR��`w�=	�5?�?�J>��F?�h?�K>{h�>�M=QL�>��=��V=�>��6D�>�:}�d�>i�������03�;#i�G��>�%?h��?���>O=þ�!Z?�&F��M��<���k'?\�μP0�>[?\��K��9���:���p��>��?�Ag��V �w�3�A�>x��<�[?WTҾz23=+�x>L���۞�>�>ὂ�>5�K�5R#=�=�g7��9��֩�<����o�ٗ潔[Z?�JL��P�����>	���ྛ�9�W��?�Fý� ?�(>�c=
B�>��>�P�r]2��]��@i>QJQ�����o�T��<���>R�ܾe�>J,$?�{,��cJ���[����<�����B�fh�FF>.�6��Q	�D,�=G(?SR.>�%6����>�0�?%���NUo�H"�>��>S%��̳%����940> ���1��>z�"?ɝ?�<n>z����>bE�=�]>K\?��t�>�X?�=$?��4?�)?Y �>q,����?��>Ԧ��o�s/��R�eU0��~g������>���u���>Ť�>�B���о����-9�<E�����g�>	5��@���V�>�)(����>��?���^`=�����-?����K��U�����^����!=�*�=�����%���н��.��ˢ��j�=Py�?|×?���=p����&=�w0?󻞾�@_��.F?��|�&`�>��=n⾘,z?Z�����ԋ�t\V=�`���Ȼ	������>��>z?ҽ����G+?�?^�8��Qn��Oe]=]�N���6��>#]�>V ?���>T%>}�+�]J>��h>�>�>
Ƕ>;{��p6�ض�>�A�?������=�?�>�p>i�Hdk>�վ�9d>�M�p����G7�9嵾hg?�i��Jч���y=*T����W�K?c�ݾ:�߼q�>��f�h¸>3p>I?>c� �.g���d��JH�Ys�>��.>13Q>��>���r�>��޼d�T�$ژ�4?���kп7�l;�Tj?Ln�?#&��.?�2`��3>i��>��?���B�A�F(�ћ��\?ƳP>�k�?��"�Z�A�YIK��M���.�����#̔�DAT?p�e?�"��u��=2<�Q����4J��ƀ��dR��+F������{<����A?�����W�>X�?A��=��<���,?��@?G��w�?Q^?�a���"����>TL�=��?�$�>�bg?�s����<��>����+�#
^����>,�9�&�����Ϗ�>ka?72>�>?(YY�ފ�=��>��>�?5���5�ؾ�A�>z���r>��*���b?Bl"��V<��^]>�ή�Y��{�H���+?O[ �6���� >�?O?�d�\�?�>[��>��;>a�>E��>�������i�>I��):?J �Lف��;����Լݖ��uʏ�Z���� ?�e���?��,?<G�>�.�M��;��b��|�?J{=�?�?��=>�T��:P�:�`��n�>�G�=G.���o.��h�>b�*��t�'�"�@�^d��2߄���?�J�?US%?@��0r�>�}�?��v?7��'n2?Kn?�%��(T?�*�>�n�?�4B>�?r>?�+�����Ɏ>;�g��k6>o����!������ݾ6�`?�ژ��8��=þQ��?�\��Kþa�l?�������?��n�
���}��Mپ?��>[�:�Tq����=�����>F����i����Ⱦ��y����P�>���=�r���ѧ���>�M?}_���&��V�>Mj?��K?��/��ھ5�Ծ9
��hM�E�D�] �" �
-@�i���6ɾ�V��F_?-�?�ľƸ�>� �tv�>��>W~�>��?�s&�	�/��F�>=[�>��\��?w�1?���=B�>L�;�h�>,H����>ī۾�p���7�@8?��$?���>P�?(�>��>(?�WY���@�bHQ?ʧS��qQ��I���!�u����J?�0r?�6�F/��ЄP8�x�>���>*���\;��J=��C>��*?^ẾT
>��>Y��>�N!?�Fֽ�7�>��=���=���<?l:?ZM�Ø�>����0"P?_ݾ�"�>�;!?m����Կ�vw?��8?�\�>/§���پa�&>�R-<2A�L-��k�x�k��>T{� ��Bl{��7�uNY=TҲ>H-���.?l���Y��>��i��~>H��>,��?iB�><d�>>sS?:">zF�>����),���?]?��q��~̽֩Ľ.e�<�Q�>��9>絷>�R��c��?
��>��W?#j�>��(?U|)�oOo>Y��U;	�3�?�W1��El>ۉ�=4B��#ڽF>cdu�����������>�y?���=�3�i�>�v�?R|�>#�Z>�@�>qm�>h ս�S�>���=��>\h��.R>�>�>�;�>4.�J<$<�𼔆�>�:G?��?�~�>��=����nJ?T�)�	�&����>
����H?'O��T���Xw=h�J�ֿ>^�_>�*
?wFe�P;�@ڽ�3�>�~��o�G?X U<�p ?��^���P�i?�$���Ͼ�m����M�M��>Yӗ�YB���]��^]�l: ?}zžYyܼ��>O�>�э?unR>E�;��[��|z���>�^��E��>�����XBi��#�>I��>I[v?���>8�侊�
�y|?�$U?Ҙ(?�>O�_��Fi���~����>PՏ>����[1>��%�`�-�>t�}>m�ʾ��?��>��>▕=J����2��6پ�~�5�?��9���B�ݪ¼g���v��`���y���5v=�_E�o��b��VԾ�U���7?hT@<��>yq�~%.?l��ۈ>v/�=\�>a�Ѿ�CJ���G�m?f>0qB>�C�>��n?��?��Í>�[]��g]>�.�TB����s>�G?#3��T�|��Y-��J~�^��>m�־����h�1������� ��S�������u?j�q�>�蜾9��>��Ⱦ���>w�=��h>ϕ��޺�>.����K?�"�>@;�? �?}@?�|&>�Y>W�8>pXE?�ǀ��8����2����?�,N?+�X�;O�><3?=3>�󖾬��>���>���>��f��5����=|��>�/x���>|���⚽vc?[<r?��f>��`<���>�o+?FK�>Ű�=H3>��>:�=����M�>@ ?DPG���:�𖾄�6��k�=�l����`�-ޖ>���qA�>��?��x�ܾ�����"?|�ྈV���C�O���Ⓙ&��>�ʾ���<���='��_YY�K�N>'ۙ����>���>��?u�J�
�s?vz��!?K����㾼ɹ���K���9�?4�B� �Ѽ�����N��0 ���e��2!�C2>���U���}�?ad�]��1?r�>����>��>��̾� ��ֆ��')���H�h�=y�?T�L@+����=��>gǎ>���0 >�=:?=0�>k��BE�ϗ[>S�><�r���H>�l~>��<�Y>�׷>�p��a�}?�@Ⱦ�p?�G��
�3�C����ݵ��}J?�2M=��8�����ｸ>h?�V¾�+��啛>�T��Xb ����>��c��~پΐB���Ѿn>��O��1��C	}�UwN���?�a�=��>�߿�Н>� ��y�H�r?5N�>@�<X���� �8Q>Gq����=�!>2�Ǿ�Y�)�;�v�>���`x
?�Jo���>0~G����>��s?t[<?�ͣ�C����
���F?�K?fKq������ھ.<?������>��>�'��q�?"2Q>r�?�	���?��5?�@�?邋��M?�]��v?�#'�|A ��!L?l�}?���D =(p?/�彖e{�C[M�����)�#����튾T����2?@q'>�"����>���Ӕ?!8>vt�>�}?,:����>U����N�8��
=��V7���>�>�� ���}�#�K>�A>({0?��>T���˅�&�>�Ὠ��=�	~>ߌ��@�^��1��J�ν�xK��؛>��-�Z��>?@v>>Xe� ��=�w�>��N���`?`U�����=�v��0>,2V��h|>��s>�?��='d���_j>�>�d��cx����6�e>H=x�����e�>�T㾞T彍�"�?u�>F� ?Hq�߫���}�@�?��?<d,���Ҿ�e�=r\���/=�Y���!��>��>�5��^�*�>%H;�n_�����3>*I�<��K>�A�>���UJ����>6ʷ�!����6̾�T?d]o=�C�s����>%͐����j��=0>ٛ ���3��ކ�
�>���������پ�j2?�>�CP�O��H�?2h�?�
|>�x���SF?LD7�DM>��ٽ��?m��;vy��Ŀ��^����>No?Y��?�!Լ��?#g�.]@X4>�og<� M?BJP?��>�����?\����Q����n>ֲ=F�#>�7�Wq����0�v��>�J!�%�F>������H?$�<�q͒>	Nؼ��=�[��}�>r+����>H=?^��>��w�n	
@��Ӿ��?*��=�v?^R6�A�?Tę�3�K����<J�>g�C>�Ӿ5f�<��g=yw�>~�ʿK�>Á>�꠾��{>N*�q}�?�v�n��5���F?`�0��y=v0�?W-��$�y��'�?�Dݽ<�߽ҍE?|S��Z�ǿ�:r�i��ˣ�:��	`>>����,��<Me��xO?�z3?����^Ծf� ��U�͐6���?�s¾�w�>�[�?�)������?^PG?{�f?͵�?"e�7�>��;�?_
R=��Y?q/3�^i�>-5ݾxP8<�*>V:�?�?I�>����o�-?�5�?���?t�:�1���I����M?.x=>�����~{>c[�?��$?�{7?����3������?ŨI�GQ�? J���}���������V*��UE�?%z�?�*?�V/��@>�p>�D�=��#@����Dƽ5�Z�h�?��޽�P���c?�V%?�m??�(��N�>T/��[�>+�Ͻٕ	�/���q���g�=��f�?Jy�>-�= [��f�t貾��?}��Eٽa/����޿(-N?��q?ܴE����>Ԕ�>��߾V�����>\>�?�&>+:����y?=����,�J�N)-=��f���!?m��(B?u?�;Ծ����*�� �ҽ	3���X6>_����@=��>H���bQ�?�����O�>/޾�*<?��?GŸ��/�?��d�	~M�>w�>pÈ>���b�����?��ￌM ?�E�ؒ?����?V?���o?8��sk?D�>ҟ&?*7�>w7B?/:?M��N$?ݑ��������>]@��~,���>�Ny�[[�fj�?����1����5/����;��<z�@��>���>N�>�aI�N�J�>o��>{��>���?GJ�>�z?`o߾�n>%١=��@����o=���>^�{�׿$]ռ���>��Q�f�?��e?��?݁.?��q?�;�@�/�%����`>�F��O�e�u����?t4����>�o(?Q�����|����&?��a?�)6?8e�> �>���1V>�>ߴ?�T?=�:?��o�O��>�45?�bB���7��
��:�=Z>�'�>�[�=Pw�?�O��^ي>�=�>l6]���;?^�/�*j?��ھ�<4?"I4�� �;U�����=X�>���l��?ڙ�<���>��r�?FN?.��>���?�X�`�l�俅$��*?��H?���?@�>$a���s��T�>��/�>Xv��b�>*�?�̕>~:2?�%ξ�����Ub>��[��P�>�`ľWpǾ��ؾ�l=�s�>�vw>��a��B�� w���>$�]?��n>4(��q"�?L�?��>�o� ų��6���g�<m�/�l>1'��]��d���H�Q	*?�f=.�>c
 ?�t�D��U3�=R���d�1?�?�#?���>�4>�w�>6��>��۾.���S��>u���fx&?N8��];�9��o�>Ø���36����>�L'?�d	���r4���|?<,A�>�J>4����y?�����?:p�>�{����Q�������yѼ�	���@��0\���8D+?3xd��_7��뒾��>��?�t���?���[7�**�>�s6?em�<p{���\���Y|?��.>n�5�˓Ѿ	x?#�>7��>�.?Z\��۪����M�k�X�t����u?2��?��쾌À?�0>��>g:`����Q��>o%,?l��=)��?���?�_?װ�> �F=���=zV�>���TϾ�G��0k?<?4�r����d��Q����f۽�W���W>��?��?͌�cך��l�;h����N���T������?L����h�o1�9Hh?������%AZ�=�U?��$>�.\��΃�A�?��+?�V�<o�z��g���>��)��� ?�ξ b�>q������>�U�>W����ռ]F?�"�>O��?I�;�_��=e�f?�)w>�-�C�>*�]�[q��"�����z�o�1����?#�1�?�ɾ]���]����>���?-��?9{d��? ?��?�4��^����>���>��5�>�蝿��5��َ��-(��d�?���>�A�?{-M?|�S��S?L�V�y�=�=� ��Ru/?wG'���=�Hh?��>a��>���=��L�g׾s���*��Í���sN>���>�>��R?������?��Q�XQ�>����_?�����e?�^���)?�F��@&?И-�G�?g�"��;?�0#>
uԾ�о#0`?��`?4Ac����=wM=��@B��뀿��%?;��'�U��cd>#_��ҵ��>m���n�},��B��<q��?ަ�>�K? �z>�oz�2g�4(�>8B�1�k�U7?�h?����I*��UǾ�l�=��G�|�?;���z"f?ڱ���Y�'Xv�a�?.�1���Ծ_��U$7�S��ȭ?� =?���<��� ?a�<���a����d����>���6�<S꛾)U��V>'/G?���-�Ŀj�?�G2�3�پ	�f��ʢ?��="��L�c���,>��B��R?m�=2�)?!��>�ʯ���?u7�?gK?�:�=fnE?U��?i�?[>ra�>J5	?`n�>�!���m�>i��?�<]�?�����E��?�o?�>N�?�P���Ё�) �?]��Q]?<�?�.Ŀ���=R���S$<-;�UYپ���~e��G��P���Wg?��5��"�?h-�>���8j>9?��a1>��,>7cW�?���"?�>O�?;@U����>��,?TK��>�B���?5%>jjd�cpa�)�>������>��B���?g�b?��1��->B�@Q�H?D�q=��g�tS�=}��>e|�P!3?���?J�����ٚ?#�`?8gj>��˿�U?4 � ���# @W߰>�g��>b���Y����	=㋬��7h?JoC�s����������>v��PD�?�'?���> �?$b��NR?�z?>R<��]�jO����B\�	|�<�na����%��=9)���m�#C�=��>�K����*>����K?��>�4>�d?�?�6۾2ݵ���m�4B�>��?�{t�k0+�:�>�8տ��O>��u?�m/�������C���Կ�i|>r��?�E{>~����J�"�L����=�?�?���=�L?s��>��N>�s�?>C}J?ʜn=�F�$*�bݓ�݁�����%����BP?�>�(>�"o>��?�=q>=�N)>����^¾�S[���K?9>X=?���ۚ��Ԃ_��*���q��A���<R��ۅ"?��4>�q�\*1=G��= �$?���I{?��?r+��i?ș�=��A?��S�Ҙ�`$��A�����֫?U�k?�#q>֔翠���6��r���P�>��3>ӌ��Őƾ�=�왾�yǻ�P�<8��߫_=�r�>c�M���U��Kt��u��0پ��=�h�*6�>o���P�>��=�Z�?C����\?� �?�)>�9>�x��Ö^��# ?�Ց?�^g�h��=�y������a_����di�>�!I>���Vߙ��j�>�  >����d �=2q#>�^�?Q���l����P�e �?��?� E��?��OK?�ש��Ԟ;˵d>pkc?뗨?k�J�~��g^�T?��(ƕ�/@	3Ҿ��>F&a?�5?׾K��=��n>d,�A��=(">"��>� :?�;��'�`��J*?wE�^d��e��EP>yD�`h4��.���a�?0�E�G�=���>Ѡ�>0t�I�;���1��*@!�l��)?6�ˉ�������*I=���<:ڛ��m2=�^6�np��&M��Oc�a]�N�=��D=|V󻖢0��6=BL>�d=�uY>9��=7��=4�<'�B=��Խ����Wн(�.��j�����x����"w�6l��y>c��^K��4�c��<�I޽$(������vI>i{�-;k�Vu�����<}�=Pb�=�Q >E�j>M���qĸ<��R=
mD���=��T>���=������/>׈�=ly=Ŧ+��a�
�5��׽B���v�b���J���3��@8�|ӧ�����ǽ;��$p*��H;��9��W	>��#����=�:>TK�=v�>7��=1�>՞	������Pn;�pK�E~��!`��Ƚ���<ws`�N_N���`F�=D>��s=�U5=�m��[<�|(�ÿ�=c�
=�#l��ʩ��r>���>��>�3�>�d�>v����4����=��=��E��T�<O���W�=����8�'1M���p��3�䌾R�~��|4���F>��>]<>yGr>p'���_�;���ޏ�լz� �b<F�9��c���B<=�5�=���!$L=�P
��Q>n/>Y�>J>�>�r>�d��
 �=i�L�Jj�=��O�F	�>k<1>�ǋ>5$�=3F�>?�Խ����bؽ&�q�rȖ=�o7>s0V=�&��3�>�'�7>�a;#�=�k�$ Z�61D�R��/���i�����(�ཞ�����$����8����s7z�0�����~墳L��=F䋾T28��<�<X/�;g㮽�S(>�Ȓ>�X =����d��=B>�=���:݌-�OgG��w�չ���ľmY5���	�ǑH;��(����=�7�>�>'�=z!>�9>Syb>p�1=�Q��>?�=��g�P��>��>甒>1�:>`P�>�S=�GC���=[�:>a�$�ƻ�kz��j[P>t�'��)j=z����d>Y�>�x�>
�>#�>ύ#�-�l	�>l���w���A���q�>3T�=K:1>9WO>��>��~>�y�=E�v=w�>���<T� >	�-��oc>��;N�{e��GZ>�\Y��+��\j=T��>5�Ӽ(J�>9�4>��>YQ� �6>9�>Y��>�RؽkM>�V>=�>�R���~������	>�1���f��nP�i�ľ���̥=�鵽�=O�>Z2��Ӄ��,�<m��=����M6>ؒ\�*!>J�u=)��=P<>="OH�Dz�=�&>��Q=e�g��_}=H�#����^�ǃ���j˾ƾ,E��)	��&��;�>T�6>��4����=EU�=��h>1�r�r�6=Sp�<�3>'A��2���-� $;��>}*��$h�����=�D�Kr������S<����|�-�3�!��)�<*����O==6^r;�= >xe�;aV>�y>ضV>
��b�\=��]=�>q �t����C�^�*<���㏾Q[���5-��l�<���꽂<n���,p��%��=�:R�E4����=6�;��>X3�=p����PU>���=��#=��K=�����JA�2�i=j���l.=��=���<�R½�%�=ȴ�>��>I�:>�>��=��=a�o1d=�m7=
\�=�3�yM,>|=���={��=!Q�> �>S�>ݷ�>���>uR�=���ލ�Xϥ<�;ViV��'��b�<��&��$5���!����=��>��{>��>$�c>+$�4��_t>�7<�OV=����4�:~l��i6���?����ٻ���*�-U�7V���s��6������+��g5����#��,��`��
�����2��<#Ƚ=�������K)=��)���ʾ��d��ㇻr�n= �U��)�=�s=E� >��Ľ�	��[��=��>�B����|e�<Æ��&h�aػ���`��=N6��`u�=��<�+W>%٘��[�;H�=�|>����Ј���������v���)>f*��xf��pfg� 5'=��?���o�6F1�>�3=� [�� ���s>Շ���=B��=��T>o�ѽF;½�и������gi��Ta������<*�O�"p���%��6 >6�f=x��<��=��8;$&���F<RZ\>|�	��a���.>P��>F�=!��=�G>���>U�>%�>��>���>8켃�!_=o/����>t밽z��=��ӽ�t�v����<�S��<m��ҷ���/b���O>N�ɽ=5��B=�<ܽ<A�=d��<?2�=�>�=aO>�K��l���:v�<��=���5t��JnW=����J�=;��s���y�
��;��	=�z(=�J���.�=
��>�N�>��>�>��ݾ񭯾C轾�6��Z�5 ��E-��w��pG;�������i���M���I����������=^�=��=��>�I��,��R����jc>/O�ϊS�A�Ƽ4;>=G�,;�z�(>��>��T����=��=_��=rSA���!>$�>j�>�C���>�P�=�4>�u��m�_��*���a�=��=�UZ>�O>&�C>U��=S��>g�>�Z�=uR
>F̄>#7�=�W��J���`�пȽ���#�<N1�O�a��c=�w>��ɽ��u��
>W[=��y=Nz?��w3i�D�Ji^���5>�Ϗ>A�=B�<�.x>eF�>]�>¢*>mU>P�>�6>��2>;��>�Ƚ>f�>�=X���r=\%>��_;U�E��M=��=.��>�����s�=��*=��>,��\������Kg=&PM��Y�ч��9�[��`���N�=͖t=��	�+����N=�N�=����xx���&=1�Ƚ}�J�r�=����,���U��pT^��󗸵j�=��9<�s��_=��>����eT��,Ľ&�	;�����	=j�=H���h�Ի���H�������M�<Ҟ2�#B�?���5��Ġd>�'>`�P>�n>��ܼ���=�	=<��� ��=m�w>���=6a��xw>�e>qV>����E��!a��ʃ�c9���T���@����qx��!�T��@7>(6|=�� �W�����n=�A�=�+b��[����
>m{�;�����ɾ^_�խ��|���も��z8=w?ʻ��=�I<�	�=	D'�-�V>E���#&=1t%��<�=�#�=��=�A�>7�>jo=~��=h/;��>'"�h��<��	���>���=���;�t�=B>�i��(�����=�D>�X���o���<��H>���g���ћ<�b>����9gO����=�i� iǾF�[�1��yt�P֞�a5q=��;���=����ԤH��o���<W���������¾3ü�,5�Gl0�!cK�R>@���UG�M�*
>�>0�.��&L=0��>�6>ViX>�ϟ>���>'^�<��>q��;��>c�\=T��<V��= ��>�S�=��0>T�+>�+�>�N�>�o�>D��>�%�>���<s�.>"�-�`��IW�=�
^>�M�c�V��m>H��=��ȼĕ���"4�RT:�|m���ǾoD��}4<��L��]�B�9��9l��=]ٽ���a3>I��=���=X-���;�=��H>B���-��=����W	�$��;	\��7�=�R���n>� *>J=�"��_�?>8su>r�>��>hl�>��r>�,7>��N=
G�=�d	>g,��ד�Y����&>����*����k����;��1��T�m/~���Խ�w>���A�ƾ�4p=u�=
邼_qž�$�>���2����Ⱦ歷�����������޾�����^����Yѽ7WܼV4�=���=T|H�5��� W>\xG>T{�=D�&����s7��;Ň�\��H��Ī���=�h��)l�)?������<;��>����t�=YhȾ��=eM�G�=\=�>(��>.":>�<>:��>e�!<���<�"=��H>S���
����A�z�&>�����U���q[����:��.�wI	��uB�1�<�cͽ�8ԽTA����8=����&zR�,���Q>]�;��>u⫽�v�=[��>$�n�W#�|��=�c���ג��>��E?�WԻ~"U�t:`�X�?���c��U糾�f|?A�?e�"?|���k?����W?�0S��?���>o�?f�?qpG�M3�l9���i߾�#ܿ	�ؾ��?߆��c>'��<N�9=X�>��<i�=��ob?<^�>附?9?V?�O(?-�˿h�?�ě�N��>K3�?��;?��>�G����?�d�?s�?��-?��?��t?ǖ;d��=H�b�_m�� �x�:	�>pm��P���f��-�ރ��J��O�?r��?�E�JH�>X�?�ĕ�9�%?��>Е�>%~?�>�E�(gྒy�>^(� �_���X�;�����l>��.<��?�͏>� ?#r��o�������=�g����S�=��q�K�f?�7�=��5���<?�}?y�?X>�?=���F�=/�r���?`վ&6��K߾-wc?�c��m!�C�� �#=ܱ�$�����^����>��D>��;?�]����k?x*?��)?�Ї���ۼ�ƶ����![��9@��+���(?�*�>^m�=&�3?�c>����Y;>3�>��d�"?)�B?i���h7>�ls��H�>��i�_��	>�ϯ�B�E?C���'�=2א? s����A��ڼ&�>MO������ 9���?�>Ұ'�8\���f���j'�Z���ȻξQ=��$�d�=5>��Ͼxtb=��(?��E=�蒼��3�م��k��Bdy?]2�?�D�>�#@���>QF�>�)�>�_?#s�<���?9!S?CC7>q��9�ǔ���&�,pZ�����L>���P�j>t&�&{q?�&l�k >wW�>)�?k|a?���?�#?������@E�Z�V�z��cC=~��>�7??p]?�[]?E
>�s��)?�\�>_犿�pþ�?���?���>�?5��?���>W�e����??|׽!e���>��?�vr���8?����gf�?>�?�!�=>��=?׊?�˾{��>H��D�=fC$?�eR?��N?؅?a>��>������H(n>�2^�*��>�l?�@?,�<H�!?]X?/W?2�O���Ȉ�=��>e����*-�6VC>^jĽ�^��H���+�9i�"�J�C�1����B����>)O,��g>0�-�9�B>�3)�{	���>���?���.~��ݗ>gf>8�I?U^�?�	�>w�ɾC	?�">?�1��J?d�:?BTN>>��h˄��"�J~��~z¾ @e?�oX? �@6ž��>���>?>�J�>�����������>��>��j��?q*^?���>9 4?=��=7ȿ=@�>==>^F���m����[>p�Ǿ`���̿���3A���(��۰�A�>Us�>c�G?�l?m$?�*���Z�=�b?=Yr?#=�"�����6�C?��6��~�>�~��w�?�t?��G!?�DQ��á���b?��9��蟾V����$� N��]g&�sO���>��m�?1M�B�R=�$���;5�>^�?�|�罅�M;0>�lL�륋=�������jİ>Z�?7(�>[�a>"�;�f��}5�=;y��b@�!-/�s�{>z�S��[��L8�SYq>�K��ĕ=��>�n?��0?��?�B�>�K�=��n���?^]����<�H>����2���tZ̾R��>�#>�n�>$�=���׈?�K)�t��)8ż���d�@��?�<�>��Y����/`�?��F�J���;>���ƾ�ѽ�xL�%j�=��I��J����>f�%���3��y?v�>�'��6ə��X�3$W>��^���M�H��w�?vA�?�?݌ ��� ?P;�>����I��>�����2?��? ����z�
8?��3�����C�?��z?�"!>���F�?P�!?A�>�s���}��&?L@>�>����|U�>c	�>>�">���>��z�. A>��E>�#��`�a�H�E��;�⿾�O�>;1n��'�>��D>@V,�fM���>}������|����>z�G��<�1gﾍY*��c���n��P��:�=90վ���>�Ǟ�	�<#i?�1�?o�������:'>�p>�瀿>��]���x�?�G?$�^?��?˜�?!T�e��?g'�?6�5?�B�;�?|-'�dM?��>��S���?�;P?��(��͐���M�D䢿6{�>"�>���M�=5W�����?��@�����p��f{?R虿�M�?����Q�,��-?v?���>/<輔K!�y��?wܭ==>���0��������=�e>��7�Ok�>@�?@GU?S��?d�7?S3��礆�Y��<�y�c�A�e��Δ��Р�у�?�0	���=����P�ƾ����_��>�;E���N?�{����->�m�?�S��`	�xXX?v�?�j��園?�g+�"=?0p�?u&�>���l�?7'�¥?9��>��?�������=��>j->F�þ����?rV�?����/�=���>������>��
@q_��aB�?a�>FY�>�*?�
���L9>���=i���� �?U���������=>�?���?���>�G =�bE?C2?�r/�!���Sн�>u*�?����!���e��QoS?��P��y?�p@�h�?=�����?��>	�?��;>�ض?浦?���>�Z?��>��?O��>��X=���}�U;vʤ��L?W�y�����G�>cd?G>�𾝾xZ���g?$U���B����۾�R���{��*�0>��b�P�����žRb?��V�s`�)�պ�G>���?��F�ھ�<=�	�1M�+R�E0>.P����?w��3��?��>�tG?��%�k?Fs?�$���t?>G�5�H��>�E�=���>Œ��E��������?�b1��=�F�����>�j�=��6��r��~x?{ڑ?'��>���>��j>�\7�GTP?X�i?V�>�5�?q+�_��XF?��?2"?���>T(��ص�=X� �&?�?m?�=?�Բ�Ѿ�?���1�>]|�?2�N?���?�	�=�ؑ���D?��D?���8�-
�?\����!?����k��!¹>@d�?뮝�*~<�B��?�䖾P�G�_e�<��R����䧾Hq�>�/׾�l���X�e�`�w&?��b?d�?.�L�O?�4�=�����;	b=J�b�)F��9��?�A@�H���r��R�?�uh?�c���j������<p�>,�H�ahR��O��&Ƚ�־�~��r�??5���<� Hm�-1�7���N(�����)O?�-:>1�/���`�֓��h	�S�N��炿�A�?C�ּ�������>�_����?�q&����>�v�>Ht?�I(?�m+?�,�E��>�lBP?��(?(O)�Ldӿ;���>(}8?J!B?X��ȵ\��􈾃4=���?�@I?q�?q��>��p<d�6?�@>?@��f����"����>n�>(����l?�s6���=��ÿI��y���@u4=`ӄ��˙<�:�>��R���?�l��^Qe?���?�=�?$4�=���=_�X���<>��q��޾���>W(���������|��,;�̘>�@�,����?�e?�OW?;3?Nn�Ν�F?��>Z?�>ڷ�>>J"=���;3H?���>"�:�A�@��~�>V�I=٢߾��`���@���<r��>�e>�2>����OQ>ˇ_>��I>�\��xi?��V��������<�8�ӎ���*���!W��?	�>E�=e�<?M��=,m>�%�><._?&��>=Ԃ�e?Q�vѡ�΃#>,G=L�=W��	���+�?<~S?��5�'�5���P<��?;�r� 
f=����!�>����d�>�΃?+��?�>��u?ӎ?	�5=\؍?#�K?ea�������6�>��>&�����^�`ɽod���?����T� ^�>�������������i�?k�>p[X���噢?*[�>Rh>��t=����!`;m<�	?���h>�3�=t���G4��ʪྔ�����Q����>16]�����T�!��v���>퉛>@B�>��\?�U?4PP?��=��Ծ 9u?�!?-q>�̩>�|.>�̍��^��ё�=�����Q����a>M��W����y?{�/?����$�o�i@/><����>b�s?�C�>�o�>']����-?Ƥk?�7���>~�o?�Zc���} ?�69?$�m�G�U�f��>��>xyJ���ﾝ�%��W����(Ž�,[���C>!����?Yd��%�u���>-y=�=�	V?��!?`?���>�I�=\�$���?Z�=����OO��`>�-<>^�<�~?��k*>2��>��F��H�om�>����&g���>��+��\��O㾩�~���3?-�=��%�=���bD>�/?�[\?���?^�]?@�/�����7">���>q�p�� 9����e�1�0�ٽY�������k��>S�>��^���ԕ>r3=��?��x>%��>5M��ʚ">�]���4��O��RMɽ�))=ou>6xݾ�Lֽ݉׾`�	���?����E��>ƣJ��0I��$>�Yս ��=��#������2��X?��=�~ԾJ�(���ǽi�Rm�>�!�=q�9>�q��_2R?��?�F�=�?�W�>yl��u�>(�=��>c+��k����������<�0��Ǵ�CC�=g��>d�V?�q��=H�>0�Μ>$*��#
?Iŧ>��?Uf!���
�d�ܽY�T��"6��O?̿?EǾ�����2�:?�?M�����>p�[��&�']��.���$�־s:R=���ྚX��?3�d>W?N���1���?>9�=�-�>,�G?@�p�!�?��>�2[?���>?�8�>�X�����>䬞�bs<?���>�\�~�O>��?�u����yož�&=6����>���>Z��=�A޽!�'����>q^ξ̞k�\�.?���>�cS�%����y>�F:>�z>�T�=Wxw=�:d?�<����}��k.��Y=ݺ,>��E��<��c?��@�������|>�X�>�A��U>���>�6c?*�/���=��?Cq?v��<u�8?��?M��?Ud��\�����>��?bP����D�����9����=�(���f�?K�Q�Ǖ�=\18��%�=��_��@?=I��=���>�W��=&�&>���hRu>{�G>����ɆN���1��	Ⱦz:�>����)j���o�P���P>[\��r��vÌ>i !>>H�>p�<�؉>j>�r?���>B��>&����
��U�=�d>:Uн���Ʉf��f�>�Ƃ�I%{�g����7>3����)Q�W?캃�`�qY�t:y�n�s>ww�= p>�Uy>�:??��>J�伃��=(����x�>�;2���
�N� ��>7�����,��Ѐ>^�.>u�ƽ}�O���J��@�{k'��C$�Βվ�]>B��"� �h֋>%>=���0,�;��>�_Z>P����A�=|��1�]�١�S���5پ�<>B�ξ��������=��<��～��>vW�<�	?d�=����U+��H�&����\�� ��>v��=�t�"#���x]>��=wx�>3��>��>O1>T�[�"�Ӿ(%�"ڪ<ͻ��F�����>h���u�9�в���Ғ?���>��;>N��>o�?!&=�֥>��=|Lغ�TI?�G���N���QM�G�q>��g�6�?��9>7�B(_�.3K��%���T��m��S�'�"���=�۠>K��^p����
>5q�]2������T)>���Ͼ��+��FF���=�v�>��<>?,�?X�V�u>D�t?I�>�%�T�B��9E�[}d�����Rg�>�3<�8=&ҍ?�~�>ד�>��>M�>��)>��>N�>W���?�?�`u>=`�=Q,�>0�2>���j�>���>����@<����>����X�P�B">5��>~��=�i��Q�>��>��N��j��l��&�<�KҾ��ɾߖ��j(B>u��׭@��̾1��>~�=�	="�=��?�D�>k�ҽU�>����2�,��>^Y?O��`�ɾ�1��� оUš=�]?�'?��'=�h��l���b�^D?��?$1�=���>�Mؾ���>,�4?l�?Y�l����ytC�>�^�9��|�?��P>h� ?�����|������>��=I�E>�K>�l�>��h�㼇���?F\�>P���={~�>�����A�T���Ꜿ�SB��T�\����4=���~�b�o�%��>>>ԥ4�{���j���?��D����<r�[=
�q��Z�����>�IӼ�q���˂��0�<��>^/6��/N��Ɓ=H����_�>ʴ+?���=Ud�����>:��=��þ "j����>|��>�zE�m���?}	�=�?��}y���p�>D>r+}>UǾ���?��g?Qɯ��D	?+�?b`a?�	��8j��~�=W�!?����R��=˥"?u��?�q?�?�kD?+��K?H�-?�b�>�mi>n��������f*{��F��ܼ>���>f��D�>��_?�X��uW�/�?� >?�/9>'�f=!���	ľ��$��I���p?=g?�hd?�!�>:/?�]a?#�:?�o/?��	?ݑ!?�� ?�Y�>*I?O��?�p�>��;���Ӿx�ʻ�u�=q
?4.ϾM�^>q�3?���>���*�>&S<?R�$?�����
���>T t=s���mw��+G�Eo����ͤ�>:?0�Ǿv?+��׿<՗=q�l>��ܾ��d��������\�=C�>C��>�����>�ך����><�=5˒=<W�>��>B��7PﾨEv��˧>*���$w>���=f�k�#*A����s�ľ²� 9?���O���Z�>�#��.?�\t>|�f?�"޼�?����*>1��>ќ׾`Ƅ?(S4?<�ؾ4- ���?u<?DH ��/>So�>H�==/�~���u1��Tp?$'�>u�`�)�
>r�8? '�>�	4���׽�+?M�M���H�h��>�_�>*���{��{��? >�V#�Lï?��,�M���C>�X�>��.��脽���>֮�?~z`�����{�>W<�>V���i>Mt���	�ux:>9���Y�cΌ��)����|z��?}뽒U��B8�_ా�>=����KQ=@!�;���>�'>��<o�?��o��tL>�#h��>�����)���i>Kb�����䙽R8���z�gO-��,�� >|<�>�6�����>�i�>^=G?��p�!]y��o�s���^Ty=�Ծ<�о�I�;��k�D�,��/?�X���K�S�^=[�x>�ż��>d	}>+��=�H�=i�9=C�N�F����n ?X�{�Db󾫵
?v�>qs�=��"�� ��=�%>�2?�=C��>�z����>��=ꥫ�w{�>��q?4���*g�0��>P�K?�᣾�R��@������Y2���	����=�h;���K^L?L�>|��>y3C>Y�0>ޑ>�r�=�l>��=?�t>�K�>t-?��cų>����/'켞���Ѻ=׎�Xz����?��m��o-���\�c�;=�?<�k?r�_?�)?���>�?��?�I?���<v��>rɆ<�����Z�=�VV>%����;��;�>PѾ+q
�2h콯i�>��X>i�>�L��}>�??��b��䋾/&t?�X��Ig=y�{��Ⱦ/�>�����>D$��b7>K�t���=�0�<��>wwc?^�<��x<\�n����>���=-|��? �=4$>ѷ����]�8�w���޾%U?g��V�+�K�< �!>�� �r]����?k]�>b�Ӿ�v=����>�1b?��>\�D>5ow������>P��<��>,�s�D��>��O>��{>�)�Z�>u`�\�K�l\A���>��<�E��u�j�K6Z>L�0�9x�� �P�>E$�E�p�;�?<.>���P�(���?V���Ƕ�V�u?F9����?�J���v?��@�Qǿ�D�>Y;v?�N��A?�{R�ƫ彲+>I$z>�S4?�
 @�d��P��-��>�=�k�_fH�F>n��@�ѾR� >ՋF?=�Ϙ(?08�>ǽa����){�>�����W��S�5X	������->c�?���>h�1>?5n?���?��t?�T���)?mΖ�����,d=���>ia���������1cd>��D��UW?M��?+��>
�Z>�k>��H�>,S�=m���C����)���T���-�.���"�>�N׾�x�=�?�_?�&t?n��?�L?���>+?N��?��������">`�`?��>+׏>���*����+�����n~���	|�Sf#>�W?�`��Ⱦ3��>JS(���`��X2?=Z"��'������Z��?���=�n�?N�?^���᾽Ī	�^%����ؾ|�ȽV���'?��տ%�><c?fK|�m`�h����>k�=MB!�ޱ���L8������O�L"�?s��(>�Z>x}��pW��"��.�?���B�;>�tP�d$��r)�S5?Lz���п������?���Yp>>��>�Ţ?�n�?O+�V�?o/Q��l
?͒�=�.��,}6��bH?��V>((����F?$�T�'��>�^�?:�M�ǺM?�'?��9�Z&�c� ��(��U�P�Mc��2?k"�	��>��">�,Y?�~r�xB���>�U��?J�?�c�?�|G����=%�?��_�%�?���>����H�>����l�����{?�'���M�7�?1�p�cwĿS�}��7�]i�=(�H>q\�>�?㿖�Ǿ�RI��ѧ?G�=ǎD?�-��i�V?�V@���?}J�?��V>	A
?1��>��Z>���I�6?GL=���wa�� g?
@X��=�i`<@=g?��S�=���Q�Ь6�L�?ֹ?��A?���>�¾�N$?�d����댁��u?����~�]�>�|�?B��>�?^?�c?DH?~���/�9`�z?��i?J�?D�@F�@-��t�0?�����>E�t�Rjr>��Ђ��� ?�:�?�Wh?��>�oƾ2�?a>ԐJ��0)�I}���p�>���+k��g�>9��>GZ�=�澯���>�?咿�R9�\)x��.��T=��?x��?)�?�O���TS���?�'�?�>�?Xo�?%�d�*����gP�F���#��?HQ?�W�?�v�?]-����5'P��B�>L׾�:ƾ��ݾ't�?�~�?z2?K�žޠ��p >Eњ��<މz>�n ?G�-��l�>b8�`�?�>8�'��=��B�_5^?;�X����>c��_3���
�=������?`,?�(?�B?��A?��>�O�=ȵ�>:��_��Wb{?�0>P��>}l��?��Ⱦ�in�>�׿ۇ����3��؅?y��>>�?=�h�>0�>��2?� þ͈J�6���t���8ž�9I>�	�?��+?�T��{�H?0 ��S�>闣��)��$g�萎�U�^>rU$��J�><�>a"?严?20�=��>f*&?�
?��>����{%?��C?-$Z�����?�������?��[?�D���kp����>$��>M%A�����M���nz=�k5?5��>�xY��J���:o��/�Z���^ʄ?Ƽ�?�P?��A>��<�"�#�ס>�dG?"�@�J?|P���3:�Mݨ�L`�?>u%?�[F����o|߿�mX�5C�&�>�^N]��0��������?�޿-��>���ܞC?(�hE�����"�@Y�?��>��	?&�>K�O�_k�ͫ�?u�(?AO�?��?�����>W��?Dkp?1M0?��,��G0��C����޿��Z?ۿh?��~?�r>r��>^2<U֒>`�"�7����9�=>x�?_�?��ȯ?��?��þV.�>)Ɩ>�p��x�>{E�?��I�f<��!��j�2�R� >�^��񍕿��C�v��҆�@S����Kn?対`�?(yY?w9.�Z�7�mYE�L,B�Z�>񲳾�F�9��4.?����[L��D��?�#R������$����k?�v�?_h��-��?�$���Ὢ�T��?�f%@8�0?��x?َ�>��P�}Ͼe��>���?P�D?:��?�EO?�>k�>�:>��?>2M��Q���{�
����ٝ?�O?��!�>����O�>t�f>��?��?�H@?��z��K?4)��$o���;��D~?�ɪ��\*��l?�^��^S����0=��:�r3���'?*h?oǚ��ǿ����A�>�ڞ?��?l�9?Q���,��� [�;��	$�?X	�>ۄA>k|Y?A����L?�/X?s��+��hʕ��3
?٪5>j�[Ky?oP��6�>G�!> �u?ăi����?���=������^B?St��'��=���>��>��0<�>k�=��4?s�?|�l?&dJ?aU?~�ۿ)�ſ�a��9>E^3?T#�=̱i���p�yջ��O$��\��Mv߾�=�?F�?�@7Q�?[<�=T ??�d�?|bX����s
������������=E�?��v�>��>
��?�:�\*\?s��>|f�?{�h?�e,�We?Tv>6O#?�c�$��=PKl��_>Y��|�9?�+�?� �>���?
=������>-�]?xa?��?�=?m	�?���=Ì?W0?�{�l?�>a&N�$����z�>E������oꈿ7�?����J
?�+�>�>y��K�E�O���X{��?���.g�<:���5�̺Ƚ}a�?]<�>,�L>%r�>v�?��e���i��Q?�Uݾ1B{?}g�?��=�`�)ӱ?���>e=�?���?�>������߿}�/���5�J�)?���>|
�m�S�����	?�o�?b�?��?	BȾn-�?Gh?�D���V9?��?�=��1�>���2q�<�m�?�}4�bj�>��8­��՟?Vy	?z7>H��E\r?��t���:��@���ɾ�l��>k��!��?��?��?ׇ4>K�>�����2?:�i��?�\�=�T?�vѾd��>(�>g��>��C�J�>"b������U��퐇��/K>}�}?������R9?�"�?'tD�Mނ>�\�[�">< ��'��=MQ�����U�?�I��7f��5>n}>���?�y��#�?�7�90�?�?K�M��=z��=��?��>�
'�NM��M����=�D?��=����p��b����=�D=}?���H=?&bJ�g�?ş�=��$>fB�x�����Z�Rp?���>z{��5��>�d�z{о�c�o�~?/J�AG�X�K?�:�>͋?C��YF>0�=P�c>eŊ�0��zZn?��K>E|?�Y��=焿���,ƕ>�"O�lp>�b�<���㌥?�9�?Hw�$���$9X?��n=�9}>ǂ~����P��>�2�{MG�ƚ�?Z�>
�:�=�d?��?��d���G?*i0�cH��ٿ�9?�?]�>)��=��$�Z�?&����ͳ�?G�����^>�??+g�Բ�?x0�>��>����A����o>�P�떱��]?=�?^<'���?�;�?fj�?�C?ύ�K7?��?���W���6ξ@����N �#�?����4(�?2��>Z�[?:i�?9~f��!��\��>bܿH徎��?��پ�b_�n� ?�u�>���먷>�nU>�I����!?���i}�c����f��=i�>1���J�?p�G�)��>�
��Gpa?v�����w�.ec�����j"�?|�i?��?�a�B���(�9?��?%����m���8N�a�w���<{�1?LU����>��1�{��?�Y?+*�>�i��Y�?CD���/@#M?c 
?`�>�e�?��.�h��=��%�����W�ľ.���?`�0}?J�\��ej��[}�yn��1ӿ^~>=�����c?fƮ�Ʊ������z��&���t��w�*�.?��ܾ�r�G�J�|sU>E=���=��#=b3&�*p>���z;>��=����_$K�,�p��KN����<�<d�ý0�>_�|;/��>��$>y̏���I>�;>k��T�q>������νf\>�ى�fĊ�3������^����4����?�> 3��q%���|=�tq>W�޽@c��nf�_ˁ>�P�>���>HJ>���>�ե�K�>>:��N뎾6�4�� �= �S��2��de>XW<=�a=�M~�iK����/�6j��>㨾���@�z�c,�=c�o(Ž�xv���=�CY=.�q�P�>p*��N��>.VS�NΘ=��>[ս_>���=飾;?#f>�?�={ܽ��K��/�=�'��4����6���6���/>��;}�ڽ�b>OZr��&=��W�ȭ�=�/
>��w��m���"0>"F��הh=�u��У/�� �>d��>>E�>�6�>�f8>|�Žm�T>��e>�\��3� ���r >>�C<�	��>2��[m�=����jžq^`�:頾#}�>�d=_�%>��#>4 *=���;1sg��6=숑�$��F��2ؽ٪Z�۱%�%H�^�ɼI^p>���=���=Q��=�I��y�=���Z�s>E��=ӷq����<IT�=̹�"� >�6:=���'X����nH�[�1��T���������<�\i�+�C>J}o��8(>]���@�G�h=�-5��jU���ܾS�
}��:;پA4q�.���n����T�>Nw��+�r>���ٔ� ,|>� C=�޽��;�7��_)�=	�����=p��=��`���p��9<R��=3a+=9��<�%̾[��|�B�� ��G��$������k%�;w/>t��
������=��>�$>ۢJ�]�=
�t��MR<�D�gZ�>6�{>!=�=vnG>�΂>�4��{=H�=Y��>/
��Q�<e���]1>Jc�=�9��%<�5P>�0�=�9>�"�>U�$>U���*	R>�Ǣ> ���=і�U&�>�~�=��D�[���>#�
>	P�=z�>��>�B9>���E�=kԢ>�EǼx���a!��->��X�l��<C�w<�>��>N.�>M�-�H�>����%9�c�>ʻj>�5���$>B�9;S��<T
�f�I�3������������P�*q�k���Fa��V!����>�I�=Z�y���>o��'�>Kz���g����>�>X
'�P��>{K�=����r�>�F��ϭ���{��3���,�ر�=���<_��,�����v�پ���Ic�>Tʡ����>�4���;��y�>;�>�}����=4S|=�xa>�ֹ���l��������y�g>I{m����={��>��=�"	���>���>�6��DN���Z��D�>!qK=�d�=��=�X>#0g>����a�=���>:�\��>*���>Mq,=r!X��'U��&{>�C��:xe�a�0���O��s�=��%���>$�>�X��O����Ľ�b$>��ڽѤ̽�bٽ�r#��2B>�$>�Q>}k>�J���G>��;��=�>8�*�_�<���=QN��6�>�<�	�Cr�>��>x��>�e�>t����'>�k@����=O> v5�����q2>�!��<>�ه<��t���>���>�>�>o�>{�=֕����	;�n�>,�����f�=�ai>�l��`7�9B��̽��>��>�F�>��>c�<:��n��=�O<�=Ͻ�y=�3�=�n���>�� �iq����&��I;b������C	�����g��������]e�=�i��=��_�ã��T�=�Ps��]��%�>:%>yi^�����!�> �<���->e���hQ�﯌>�3=|�H�G>[��x��= 1A>���'����˥����C�=��-��I�=5�J�ns��<{>�P!=�7.�o�:�#���?=��=C���徖4ξ��׾<_�=������g=�)�=ؤ><�q��a�=r��z��>� M���;��vͻ��?�i�=Tt=�5�>���8#��U?c<��=n|!>ǳ}�N��0<)�=y?��[A�q&��f��>�>�N}>)�>:)&�D��1��$~>���Z#��3<p�,>x���d��[7��<��=l��>x�>���>L�>�.�>~�~�:d>�+��uz ��Y>��=��g�]	�=^
�f"�<��i>Ң���;�a������������v��;ڂ=��/>��@.2>	�@���߽�	S>��=��^=50`>F�H��B!>�/�>#꥾�i>��2��y�meA>L�_�J��y۽��n�i�=��=�Ka����>v�>�ɨ>^�?A�������������?0�@�'���>9��Ju��U�=jL ��uY�TĪ>�l>��#>����0q>i
�=�t=�#�>��>z!ƽԖ)�&��>�l���>Ľ$����>A�2=����>LN=�W>��@�8�2>U�r����=��{�e(�=$��=Qw�=e�C���Z��ǆ=t>7w�Yg��^���ű�o��>X���\|�>-�>7<ս�ń>��o>B>ELW>�X==F��>�^���,f���������㷽#r�>T�g=6[����6>5�=>p*���Ⱦ��=>1>>t⎾��C��+j�f�p�lR��L���+s=^_.>��0>?��>x�?�#*??[�>[ +=�R�>!3�>�=�>�J?4��>� ?��>`Rr�<�>�^<��>��������>�ue>�m��j�=^�=�S>Ӵ���C�;��IM�M�b����%[\�����R�<��=�q�?�>$!C=�K>p��<GrĽ!��=xX��[L۽*�
�����c1������f7>��Խ/�>����&�2�=D͓�[�r=>�=a�����:�*>��&f�=��U��:6=�RG>3���-��p����?.=5�[�ӧ����>ɸ?��?�2�>J�f��j> DG���������>�ʸ�Z�w�I�=������>m�=���N�PI߼�=�k��l넾Jj̽W‾}ʾ�1 �*�=x[��ܒ� %R>��=��7>Sx������>>�I=Xe1���I��wż&�ּL�,��#��q��>F|���>�hv��x�=K�>�kL>@��!��9r�X=f��=��g>�f�<73�=鹆=�ٽϘ=�u���=>��<��8�De����=]W��Ǻ7>1]�<�ѽq�^�YG�>&�����x>�(��$�'�^a�>�C`>8�得�Q=Mؼ�z�=v>˾6嘾���ZM��h�d��g>Ԏ[��>(>P�Ǿq��[��>��P>u֬�4��=��<�K�=@�
��̀��.���[�/����="��sbμ@��=C�X� ������=K]��p�>�r
�2T޽sC�>d�>���>}��>w^=l�x=~`A���j>Q��=� �s��=��l>1]�����<�
�=���=?_�>���>a�>qZ�>�`ͽ5��>���=�a�0�>��b>��;���u�;�o�<h��>�	Ӿ��M�K�S��#��-�u���&�_<��a�K!��"����i>��<��=�>�T��&�>H��=@<彶��=��M��������W=�3+��<�6�=�f��Ҡk���ýP�0���=�ػ�n���3�>y�>k�g>g�>��>�ږ>k�>�bC>���=�{K�o�=c��=,�>�^��VNS�r���M�>�3=O8�Eׄ=�E<���=���K�־~g>,��[R`���ܾ���A����=t8�F罾Kꭾ}�V�4����m��I=��@��O>/�=*�=����>t7>rH>�#�=�����LK�h�2��:�=��l�m����x������4��,��>3�2;�Lf=MӢ���>>cE>�]>�p}���=\��=��_=��>[�>��=,	>�u�>,J>�l�=��=x�p>sjw�,��<�����?S>�=����>��ܾl̃�ٗ=�(���L=�6���i>�J��%a�;i�2�(�N��E��"�>�8�
"N�2�>q��=��4?
�� ��3�#������>6~��������=j��r?��&?HVܿAZ�N�־���=t"c?��C?y�>u��=����3�^A�>������0?�D�?(��܏�� a�J�|��鍾b�#�](>m�)�%�>�I��{i�?���`)��FU���t�x'�I��>�q?�J&>=$t?�������oM_��fQ?m��z^���g��	�<���9ң?��f�Ӭ�= ;ʾ˚����]�7�=�����mw���O'����Q�SU[�3�=�*j>9#(�K��-�?�#7? =�5(:x�?�nQ>6����3��ʾ˘>]	�?�I�����Ю��.�>�4�����t��H�>|�>[ԧ�	�?��N?�S�|x����]�a��PAz���%���D��޿=����׼���>z{�=�3q?w�N?��>k�>^�C��	̿�̣���>����B��Y
���?��%������<?b���)�����X�!M?��?�3>���;�L���q?�K?�`m�}{"� �����FV�!C�� �ߦ�>�wӽ�?���=��?(����z���K����B�>�w��E꽎0�F�ÿ���>����u��A���"G�>�"�>$�;�;��?G�t��:)>�|�?��0K:>[�S�Y�>@����F+?x�>h]^�C�?�)vh?����j9���C�p�����5戼5`�?	π?:V�?&識
���=���>�N>�6�>~�=5�����?|'�>���<.�;?m�;?A��>�&L?o�>f����]��ýp~���%��X����̽��о����O��=��#>���>1�?h�0>KQ�'w����]>x"�2��?K���A>E�����>%+�pl�?>j�>��>�Ek?R%W��ܿ��9>ɡ��jC=ٕ�>Dj�>L�ڬA��
?W������t���y�M>�����?lyܾ���>��[���ؽ��W?�}:?l��h �>f2�=��?0�;>�P?fXd?5T@?�g���>2�T�\u#?��s� 6�?6���q>u ��'��<��(?aA\���'����>�}�.8�=o���$
l?&'����>��꾧�>$��>�g�?�(��&�}�m[��.1���V�<���*����>�'����D�n)*?�2��x�=X��;�?I��>��Z�I�6?s�>H�>��8?j�>�,}?�� >썊?�d�C34?��>*�v�?YI��@+��P�>�hb�%�����Vy$��إ�_z�?\5
?R��N
r�� p>v��>>�?޾��=�(�?�#�>��Q��D>�3F�s�'��#��>5V?������f��\�>�.T>t��>��1>^���d�������$?@��v��>���j��>�	L?�Mн�P?#�<Q�˾D@x�\���e?>%F��t���"���A(�:�侣�C:��7?4n;? �<s4�����\`C?|X?�f�>���?�x�>h���5?�ޱ����>��>%�����c>��?Ҕ��Ӿ�ԕ>փn>��GGM>񉠿����� �>��?�)X?�a.?!?��>+? �>����}��<
,��lO=7
����>.�<�T�?v�B�}����Ծ�� >�:V?U/-?�\�?�i5����:!�XӚ�"�'=x�g?�%?n�?עk�����Su��V�O��>��Q=ʘh? Jw?�.Ŀd:>�i�?ܸ����Y>-?��>�Q?��H>���
�����V��S?�93��i?���}����m)��P��0?�MA�󇛿�7�>�?��f�qD�!�����-�,!���/9?1����E��[r�?��?r�'>!�?�_�?\��?ѡ(?FS�L3�?�Q�?�[d?.��>䲾��+���øi��{�?�#���h�>f&�?	D>�]?�DD?�0��IL�?�wͿo�>*	��b�/��ս[���f7�����D���c	1��;?���=]����0�I4�<a=Z��Wh�����>�T�>h�?HS� G>Z�J>4�o����&{q>�f8>?9Ǿ	/���h��u|���n������x���>�<���q���.>F�����(���^�=�\ľ��
�� �z��>h�?�F���8�t�KH/>-�=��?w��>��?`�i?'�
?�_����?z�m? ߲>37?�-T?.l�>�k�?�X�?"�>eT�+ꕿ�����B���l>�;@:�μ 27>�>}���H�l��=�H�?���>4G?���>ǧc�Ya�>��?���?C��>;��mfa>�:��Ѻ��C���O��.���kF?��?��@?���8T����?�*?���>�А?�2|��Dy���>�x����>�����W=��}�`8��8����*�{���='��D['�w��$ҿ��"��˾{�?��w�+�>ߨ=�y�j���n�<�
�3�>�ls>��0�Ly9�2>`F?���|�}��V?���>P�¿�B�?x(�>x�^e�>u���;�>ʈM?D�d�ז0������>�rD?F̥=�`;��B��>�o`> ?6 ���h?&˔?Ь?�i>?*O=���b�'��
�:����<LS
�J��>�8*�ɡ=�B�?�@�>���!Cz���?\�=>[}���俽�2?���Z�P�4;�=߼~?��Q>�Dp����?�/w?�q?�j7=���?�?]��>K�q�[�}?�i?�r{�'�I��d �&��>썯?�ν-]����A&?��*?��W���n���>�J�?�֒���d�o"�Lz�1>���J׼��]p�%��'�?I�?�z�>eL.>�a	?�Վ>Ҁ���'c�y�=pF�>�j�U�_?-��x祾N��?F���nK�>T��T�=;p�7}F�C�@���>F7־a�?���������"����C�>���>�A�;Q��R?ȱ>g�Q�+����7���?~j�?���?;E?L=�?B���n+�����mM
?��,�6�>��V���?QyY�T��?y�����muR<��/� �@��T�?��s<r����w˿ߘ��B~���u�?�}5��?E�?�L��6>"GT?!�.�N'�>_�!?�2��W	���OS?�WS>V"���,�?/ok?\�6��~¿��'?T֏>�?��˿�ؕ?=�U?D�a?$�R��>x+j�X��q����>S�>v��h��>I�޽ Rm�ޭ�?v��>?�����o��U>��Z?�T�XSɾ,|]?��M���D?_?@�O?����;��>��Z?}�Y�v�r�1G=����>:�ɾ�ۆ�W����>zT�j#L>���q��?ΌP��璿 �/>�~�?>o�Շ�Q.R>/TR���>����B�J�s�9[�? �	�c"�>󅳿�Z�]r>���2�=���$Ȓ?~_�����jb?�>�� D?��G?���?�>�e�������?U*��7m=���>��˿��?Cm;? mj�� e?K���)TU?
���(�?���>����A��>ؼ��>@��>����uH���ٽBð������<w�!S�����Mt�� �BZ�����>G�>	M#�~q�?�=ufL?��>�n7?�G?��3��ߛ����>�j? 놿�d���> �??GǦ=�~�>�M��;�ƽg= �MO?�9�?�1B?��>�Y?�5(�@���Qg(�^:><���}W��X���1�T-���`�þ�fL��`2?x�v>p�K�1Q�>��>�.#�&]��
�.<�=���h��vO��6WC?ʠ}�Z���>�2�N:徏�'���c?�y��n�o?����쏺�rn�gܺ?���>~D�k�*?�j��{s�><���V��>{AD��-8�`!���� =A�a������j>(?o�?�%�>N�>e�|>�K�ϟ��BL�>��(>�A?�N?��?qV9?��>/��?m?���>z?Ś�>6^L���B��jQ=Z�?�I�?;�<�iΩ�@�T��7��0��<��N�SL�Eu߿٢#�'쾂$��P ��6���>?��뾺�H��:��VIU=�f?Ѷ\�))��`s���d?�a>t7�>������ųF?���>���>��,?M?�9^>�)H?SV?��tE��s���6>��?0�վ�%�=�O�>t�4?��Q���?Ծ~�o�A��n�����-�>k@�K �>��*?�p��Q �=z�Q?S�a�*�����>:��?扙>c�!>�?�l�>[]���	�?����2?�����]?����_k?p���;�>�}�Y�?7�;>S�;?�� ?mnX?�hþU>����������=�X?yݔ?���?�Ʉ�]� <��g��k����>��g�ڏ�=�w�<��?���>�1�>���=��>r₿�����O�-�-&;�W@�=�B�0�`�ѵt>clžU�ļ@�Y���?Ʊ?�� ��j�S���.�>+����������>\����\�y�>Y�?�W?��l>�?�ؿ���?0��ڑ%?si�����>=�g��K?� ��5��=�>���.�Z=��]?�ɘ���K?�T�?��?�>�F
?��ƿMS��>S�����:37��OL�.�?��X?�2^>�p���C�=�)�#g�?(C��K��Ɏ���i�P� ?P�?���?ڠ�=)���*Ş=��?tʢ����8x?�x?��>1���(�w?�RѾ���pn�䤃�*�-?y=>v��� ?X��>�6�Y�Q?"T���������NCο\�X�TL����@��?tvB�C�?��=iA��/ ��t��%�[?�t�?��>ᔥ?�9=���#�mҁ?�K��\v����=�i�>�>�� >�K4�?l�>�#?�|�'�>ғI�kꈾ����d	��lED�Y7�8Ì?�˽��R�?�����ʹ�΍���D�'�s?C�O�1^��n�6�2Q���E ?B����!?�
5?�%?c����<�ɚr��^��D��$�6\l?�;��E��(����?�����>a��o?�I�>>�=���B��?F/??�N�?�ѿ���?�d��OvU���l��?� �>��M>L�?�?`?'W���X,?������=��e?/_�>Z*��<��>��?�Q�)��>8�	?�ٿ�]�?D�?��?�x_���>�@k\�A,ξ��4�ºm�2�B?����,���>���>]�w?P�+�ǡڿ�Ӿ�$n?���?ڧ�>�s+<C_~?x𾒜t��z�?���>ٹ?��?��O?*腿%V�?G�?ì??��a>���> Q7?E�b�y~�?H��?m{]>h���Q�����\=��:>pe����=V�?�ڰ���ҿߓ}���>���?7��>����=��>�x���?	�'����^P���t�[[m?��y�N��Aw?��K>L��9 ?>j����������?f��bA�=�Պ�}�?W0�?-�?��?tG�?{���'I�BV�����?s=��&ꬿ#�8����>�T�+���g>����ὡ?|'2?_��>�W�C�
?�R&>�En<a�޽��=˘?��>�߾���?N`�?��>��D>|fE����>Rұ=tA¾7��>1�> ����_?5�Q?f*?�P���`i?�?���>�cý^5��v����9?���?��,[<Fբ?���>�f�=�����?;[?��C?ȵ>�\��3�>ʪ>�8��=���=��~��(�yȾ��7��ZW����>ޅ?��?��?P3�??�*?
�(?l@�'��{H�S�?+����eo>������?/���a����A�N��>n�?��r���߿d��������o[����� "�?B�q�#o�>t�.� s���>�$f���%���>o�?�X/�h �?�ّ?�X?2ĉ?���>�KO?P^>'�?���?�W\���$��G꾡�4��Q���0���գ�j�ſ��?���C;���/> ��?v|Y�6@O�|�E>�I�<��>*����%�>�C(?�.>i�=�d������E8��M�p>�]�N�=�&R���K�
��<u��Ѿ�T��׌?�����_>�$>:\6?�凾���=���66
?�~��MV׿�4t��`?i�Cq��&Ѿz��?N��>���=	;˽�#��!�?�i>������=٧��Ϳ2᭾�ֲ���?�����T%?lq����s�ε��ݢ��֗?��>��G?ΰ ?3������\9�;��>9��������>�K��2���ks����p��Y�?�v�?�п�0�=��?�<�����P���>'ٜ>h�$���>w�?����;ξ�5���^>
as��.(?��7����>�M�>\l�?4�;��[�?��?nr��޿ߴ�)m��2	½�#�?�O����Ӿ���$�����?��5�Lb?p��E�~J�ǝ�?�c?�g��#m����>o�z>V�οm@?���ǻ�?�,���Ǟ<&�B����?�����$�2̾��?O�ʾo�+���#?�¶?�1<�f�@�β?�	��@��n��+�i��g#?e~!�����sc�=�꘿���U¾vxl��	>|�g?0�>-�?��	>��>F�ﾞ
?H��?k��>S֙�������þ�l�P�"��>p��N��>}��ٖ*?��Js�?�ai>�!?�XȾ�7�? ���w?�|꾻达#�,?��\�\�?"��>�?����kV���?]?�ܾج����f?B�h���>f��"/L?[�>��>��z>�0Ҿ��@�m/�b����T���?���=��>޶9���
�D>�Ƿ�x`Z�����<�#>�x"�];�(=����>踽�>H?��?%�z?|#,?�?���?���?�?�_h>�/?.??��o��@���?�d�=�#�����c\��O��>��%���?��2?k�F���A��>K&�>d�=���D�Z�U:��	�p%B��e�����ʖ7�ȶ��k�5>ݎ��9?Y�@����?Ui?"�!?�75?!P�?��H>����E "���
>/�6�)X��)<�-�?-,;>v%�?��ſ6��>О��x?��>=,�Y?i��>i"��!='�w��s�>�#;��u�Q�ǽ\��؜�f�?���=��>��?��>����?��`?��\��;���w7?j�o?�}⾑9���&��0�߾Q�->/��4ce�ˠ���!����"�%� ��?�?ŕ���U�Zԋ?�ъ?�@Yu�����'���Z?M6g�6�[?G�,?�h@���׻?|(3?ia��ڏx��H���}5>�+ž9?T���P��.�>/���^g=g�
?C���F�>��?�"?ϯ��P��Ѿ�XH?K���ш?�j�?�C?�����0?		�> ha?h��iᚾ��?`�i��>��$9ſ�׷>�W�������M�ύ/�B����6���J�}/���g?���]��?l�?5����l>֗��n�׿V�>��2=J쬿
QN���J=(�>�8?"LT�ήJ?�g���>��?��=���>?���գ?N�f����?Pz���{<��J�`$��pK��������{�k]B�ՑD>I�G��@�=%U)?H�D?8�?:��?�缶���[Z���s?X?�R�Ϳx�?#y(��
���?�q�b��2�w>��>��ѿ��`�*�V����;���?Q�0*����=��7>�I
?�Y�>xV�?��>P�+��"��K{�1���a㿐���%W(>�3�9Q˾����ǻ�ns*?3�?[�I��8;?��}��['�-����"�?S��
!4����>P�?�?�����5����8���d�[�W>���M:z�kr-�٩q���i?�G�Ra?�iJ>�4���O��j?.�̿Q\\�럿#� ������B�;��>�/a�)'����@����%?�K�x"�?	PA?0�_��|:���&?]�f?��>��rk�8U?Sh�?A�ܽ����@�>�+?Ō��q�ّ���`�Yî?�T>��̾�&���??��={���m�>�k�e>D,�>M�Z�+����)Ǿ,w�?�)Ѿ�Mi>$ԾS�@���?�+���~�<�.&>{@�>�O�{p?q�»���>�2�=�X�Ӻ�(�>ex?�#�O}?�B��� ���]N?�6 ?���?�|?�<H?/��>Gӕ>�3�?H�t���>�H<?�|<l��>�v=�T>��P��N8>�>?SP������?�	��b~L?az��\�?k�=&�����^?�n^?�E?p>�ѻ>n>i?��a�������	�=�ھlk!�Bو?�A�=���=�m�>�-���ľe�C=ip�>��u�X�����ٿ^���5�#�����`��
���<��D�?Ob���?��䗗>ȟ��x�ܾ�:��x���+?�'����� =0�+�����o�����8oѾ��ÿ���FlѾJ�=۫�����<��>.5}��B�>Cf1��h ?�b=�v����>�W���>D��g+տ>��>:��?�e�?o�?���?Hn�3��o�о?]E>���� 
���Ǿ���9��%� ?8�����?e9��SɌ��Z9>�Ƕ��sX?Dm�����>�ʾ<)?\	���=Uە=��!��>@~�aW�>�AZ?������]������>�Q?&�(=~�<?k��)A+?E�>]��>�E4���a>@	�>t�v��0�>G�=P��V��?iU1��|�>1ۿq����=�5���?;&%>U�?��ܾ���?�y��oG���؛?7v�"D/?7`�f�p�YG���a���T�a�G�?JH?H�7?Q�����t��������>�����{_?,t6��Ys���=2�>�0N�;T�p�;?r팿8??+1ü��p�@ �<!/>H�n<�.?8�P���>
�?�a�>�;U>�Q�>c`?b>��:��y4��·=�w������7>��#?��F�<�2?u��?�i=�a�>𗱽���>ڨ�>�[]�A���I>i3�9��t��>�t(������Ot�e�"�?�ڃ?@�>�1�=��x?�W�?Kr>�x�?�_h>_�?�Q���$
��^}?��M?����"@�>t�
�������?R���#�Q��u	�v�N?��??�o���7>J�K� ��[�*��j�w�>�>j?���>�;X?I���f�>�R�=�\�������?u�>j�?��[�#��>!>1^S�6r۾Ǐ̿t�>��J>�n¾H�ѼEgn?s��?����W�=�\%���"?
<�f�K�M�#?>9a��֭>��h?ځӾ� �=K�.?�g�<�?����(���R>T���QP=����/6=:N���>�Mc?��?�\ƽ�-?�R?�<�k?�U?'��>�F�?�������߉=��?�?�� >��N=`�𾪜k>�x�?hv(� ���p?��?�K���w?Uv��1y4?�����b>����?~��?�?���>���?d�=?�/{�F�=CG�>9�>ӽ�=\Ҁ>LvT?x=?��>,��<�)?�-?y�#���!>�P����!���羏�A��8>�	� �A����_�>}���J�1�nWW>��/?�����?�C�>>���H�f�\s�>��V?qڊ����T?B�̾�xÿ�)b?C�>>��?�"?�x/>�\��M�@>������>"-��)>�B���r��1?����Q�>���?m-@>��=P�¾iu�=)�m�D�k�bs󾱻1�Y���k?��->Ra��L�çZ��#�=�m�>2��#�o>��T>l�>����=���\�=�tZ?^F�<�vY�����ze��B������c)?�>5�d��"K��i��=�?����@���2>o�[�3@��"2l?k替��>�ך�'B�>LGM��Ȉ�ɩ�?b,��=�??�(�?X?
�>���=�x���k��J˾�K侌�	����?�l�> �Z?M�J�8ޝ��O�T@��2���ك����?a]?�00?47��O�>E��u�?��x>u�?���?���Y�S!��q�&����=Z������NG>A'־,ق����F%>�A=')���k ��p��R��>
�<�u�i=�z+>����Q���7k���+zA�]���T��&F��0v�����#��f0��K�)�ÛD��*�G�n�o(�>ȭ�=��)��諭�s�>!���j�@>u@>�A��߸=Z� >3>4��o�3>l�=��:?���=g<�E� �#�z?�Y�=u�?��?�>
p?�?٘�?{u�;�A@�쾓���B⾵�n=|[�V��?�}>&u?�b?���?f��~��>uP=�'�<v�Q?�-�?��?��?�z�>���?��>���>AP��;>��?â�?���R>F���&�C���?ܱk?5$=?��?��>{z��n���;��i0�Л�����|`G�)4��h���|2���p �Zx��X���B���������=�?ǿ�.?o0;?�?�/��5h�>�]�>�v{=�W�?�C>���?&�1�E;f�Z�0<�77?�0���?KR?��? n)���F�?מ�:R��=��۝�>�PU?��?� >މ½��>�{>����E>�#��@W �gnM�;�̾�JS��䒽_KN�r�y��>v��>�'��cz���$�=u��5[�eD��ǘ?��>,k�[^>;;?]]�?�T=��>	4r?~�ؼq؞���ս�IM>�"A;���|=j��>#��=���I��>��?6�?�vʾ�rk?T�K?g��>ˠ?<X�=?��_>&�7��d�����*�B?�;�p��?Y*��ǜܿ c]>���>��������>�Ў=L�~�kN��*�P?�$���7��K�>���m_
�����k?\�.?���>��!=F(z?�C0?$�;#�<��S>��>�_���(?ޞ���y}?7r>�O�?�fh�8*2?��2�YH>O�Q>��@?�Z�?�!-?�!(���J?���a/��;8�8���2Mܾ���'ȾP�5>ͧ�>J�O� �Y��6пh�1>Yb>�j��5���O�?�F������~?�w��ܼ6�[��?���I��==�>7_�>H��g�)>M'��#�>��?i����>f8=�o�=�7�?���?�Z?_�3?Ҍ{=�}�>�`@S�=��8>��?��?X�>2�+�@=<�(׽8��?1�����?�/��D�>պ��Y+�>ag�>r 齆E�t�=?j�?���>�#�?�RR?,�޺�	�?x^*���?�E�>�V�
v�Xӛ>�f�?3
ƾ)lA?�{(��M�( &?�F>����G�>���?5��?}�<�-��>��=�a%>�W?+�*?��?�C>S?Y?{!���y;>�%J�J�ľ���>��?��E?�K?�,ӽ�>c-G�/�+�)��<�	?�zҾ/��l\!>���RV�?�&���D?��T?x��?�"���5�y��?u�e?���D��>�󏿯��?s���@?ף�=N,ž2�V��HL>��?���OM�Wc,>���>%����mG?�`��� ?��t>���=$舾G}7��Ѿ�?��ݾ�k��Ò�o���;m���M� B�>.n?+D{�ơ�;AD>��z>�N��2�����0M�>��A�:�/>�r?��X?�%�?:#?M�>���<ޜ(?VXk=8���(�c?Zz	>�*?ㄨ��������>��a?�W|��7>p�?n����F>�@��;;)�r>2��?�>?8�>�?���C=�~��:�'�B�H�!?+�=�eο�����2�*�Gi���I�G�������>&p����?-�̽�����>Őɽ�X�>�Y(�@����z�8���AS��J�Lv�q���L�>�+>Cn�/!)>�������>��9?���>2Y�=�1�<�HQ?'����=i��>�˦�H䠽)pY�E�"�/�lM��Ԛ���2��/�A�t��v�>)∿I�Q?��>E�J�ѣw�}��=� �?v��>�J\?����$��x>�Z�>�@W?yȿ��5��Ê>��?y�'���=ĝC?u����??i�>��f�~r��)z��2S?�����A���i�>�v?�����D� �;���?�7>�tj��W>t̾>�_̽6:!��ȿ&��>9����u��:���J?���=�Uֽ���Su'?��¾�~��¾��>JW?�C�?g4��Sʾ�P>����Lɬ=[�R?GÑ?Ҙ�?��T�.k�=�<0=�T�>W�9<�i�=*���*e���V?��N>r�.=�沿��B?�O�'�۾L�y�NDU?�0}?^�H>���>y�>t��>�5?��?.C|�ھ�#>[��?�����r�>�Me�78?�B�4��>��k��L%>�b�3�O��7Ҿ�i�&�@�=�_��y?E���9��?��Ѿѱt<ڴ��d�@��$�� ��D| �I����>����ѱ>�i�>P/�>��o��s��X>�ڞ>���N8_�>��'�?;��0�\b>��:?H�>왯����]K����?�=a?l;\��Qe>
��)*%�}rҾ��?��S?e��?U5v?"�'�	�>�(1��p?'�-=Q���)�f���|=��.�ھ���L�>R�,?��n���1?G@A?Z��><m�>b�7?�yϾ�\���k׿h��>NO@?��q�Hm
?���}�^��j?X弿�& ?����Ap��$��>.m1������!@>�\�>���>�@⿡�X?�YپY�>��?zk�� ���H��\���6��[��u��>��a?`\ξhK���p�?+�
>�����~������ۼ3`�{|Ӿ�ZG��ڜ��+>���<\�O>-ҝ?n�L��y]?T$�?1A�>�V����y��x>@%�?�>�>
��>�l?�ڠ�5e?��>a��?��`�m??�|�>]	 <KԂ�1�,����=��>�1>"F8����UV���Ƚ?l�>�:-?m�;��\�>�6u?����̐>�eԾ��(?��2��T�>5VM?�Ӌ?>Y?Te��;�j���O�n��P�>��J?�QD�����
?��=��j?�����/ �����_ɿJ��?�%x>̱l������&n?悛?W�L?�Ȱ���2?�VA�<^�=�C�>�'�?�)?���>y�?�+�>E�s� G|���X���>�x>�,
�����%>V�?d?��Y�/p3?�C�������X�@j�þ}�O�8'A�n	+?�>�Pƾ4��<K�?�I#�����I����=�������v:����E�">"�t>�䗾[V�?�P�]�徵X�=e�?�8B����oR>��9>1?��>�/�}/�H% �� �8��}��c�>�~���.�P����Z�>�V�H��> ��Լ羅�%?ܺ����?�D�����%�>�ݬ��U�<�="#?ab?
ؾ]�>_���>�g��Ts��&����>�[�=5,!�xz�(��>`d��n@��P�^��>�W�=�(V�J[6���>6^?�#?��4?E��?������c��ld�D>A�!�j�i=�ÿ��M���\��~,��v6�����B�9������>��G?�N�r�龂���L'?2���,(��l+�����?���=+���E��
�?
�j?�ƾ�����D	�d��=���>�I>S�E��}�>��� p��%4��+?�Sb>Ũ?�u?jJU?qz��bʓ��,'�%ڊ��,?z ƾ��Z�Kþه*�2YS��4<g}Q?���?I��?��?�{,>�����PV�����
�}�����k
����Zk
��]
�����1���&�?(?$�?���?rˌ?��4<��h>��h�OLW=��J�Y��=�(��Y>t;�0C5�����Ϝ�S]?��=���>ʲ@���W�Z����Kq�>U%��SK7?�%F��w�>x�>�R> 	нS�.��E�S?3����j��7��^�?��K?*,>�����%��0�?�.�>���?i��?$w?�Z8��<f=T�����J�|�H��U�>��?D�Ѽ�K3�V6������["?�=s?�kf?څ?h�? �K����ma��ٙ��3?*��r65�*7�>L��>���� ��_������>���~�����0�>M@?̂���G���=�Bl>>������T ������=���H�3?� ��d��i�i�Ĥ?��>�-?U�:���>8j��]>�@i?�/�>He�>�7;�E[Z?��`��_��!;�>��?�o?%>)?�!O?�#}>�a�ڤT>��?P��>Y{�>K�޾4
�Z�>����4�<?���?���?L�����R��of�6�B��V��>KS�?QV	>tDz��&?��?L0��K�>��T�(�>�Pv?�J-��=f�iMt?�#L?l��>|gؽ9Y��ղ���8>.�Z?�q> IL�@��>tS��23>��]�f´��\1>Ƕ>򶣽G����4r>r/��u���J�n�*=آ��R��_x迏��=���#x����@���(E?�	��F�����8X����?ޣ=�O���9�ea�?Ľ$�/>6H���?AvŽV�+�ഢ��U�?���>0���n?M�?��>��)>SX�� qt?��n�{>Ƽ���?���?����OH>�M/��J)�D<̾���=��\>.J!?��?I���S��H�>>݋>kN?�̅?���>2� U��.e�xű�Q\Ⱦ��?7��=�-^�[��ʂ,�{�u?���&p5?A_@?��$?��/��6��
x���&��/¿��>���>uĔ>����}��=�y??�b�?�Q?�*$�i�5?	o�?�Ve?��|>��>��?rT�?�D���v�>D?Ȳ�?򋧿V����<=�H`?���=2�]>f��>���?֢N���^靾b�n?������p��: �W1о�C=Nng>q?� >U�q��8�>�� ?"��=�o��=�>�>�����,���¾&�)?�M@�6>@(<��>:�?����d�;�(�'��ڵ?�"`���?�P���u?�>.��ݍ�L�����Q>ϥ?ϊǿ���O�¾�H@�'u2�0�V?1v�>R�R?��Z?��ϾeE?tnh?�f��B�V���>S��?�����_?���t��s�t����:��
y�|I��a�?�M�>��?xc���}=�/��,�=?i?7��Om�3��?��>J��>��*=��h�����<���畽���?~_@f!�7�����¹>@m��O5�;���lA~?��7������J�>�I�?>�����������{���A?��ds�%ھ�'G��Æ>Vz��0��N=��<��1��jȾCwL���վ\�����?�����H?Jk�v� ���ؽ��-�u�<?9d?fd�<dGW��E���		���K�}�"��?>��?�V���z#>��ؾ�pT����VE>02?@�?Q���\ZY����da�P�{�B��Q�i�(>��;���=Rꐿ@?�#X>F�>��">⣵=��T��K�>��3��@�������þ����)�=[��>���>��½�7O��8��~B�>}�>�C?"��=p�％�n?Ùɾ�5��P7Q?=oe?sr��|U߾Ȇ���:?\���;��?=R�?��?י�s�����E>�7�����S�?�*>��k��i+?ѳW?h�?��?8��ty=�&�?�k�>��>�W��/਺�
�?���=��K?i��]5P��rL�6v:?k�v?�"��Z#?��=��� �?~�g?�k�>� )?x�=�j?]�\?���?�<�>�z�#���B��1<�^a����
I&���%V>��w>�Q�>�/Y���>p�?�V�>\�b>�M
>�H%?@��>�Ό�o*T?|��	I ��`>c�>�l����i_�>�^�>���=%jF���=\�_?y%?K5?si�����n�?q'�>| >��l��2�>	 �>�Ң�k���f�ھT�6�`��>�0��9^ʽ�:'�"��?�i���*���?��h?����wM���>�y�>�P?�H:?C#�>3� ?�刼WM�ǃ/�lж�s�	>�G?�賿F���E?��9>��?�D�J�F?��X�yd����9�w?>��=Ō����(��c>�K�=�
�����Q?,eN��4�yR��$�ڿQ-ԾT䡿���=��?�N�å���7���K��h���9ӽR�h����h<?w�.>G��?ż���-?Y<?<ϧ>��M�f��>�X�>�|��$��>��>1i�>򰾠 >�-�>��!��U��LA�(�������=��R��\�*(0��"?�*%��a>N:���X���<>���>'?	�>��W>r���!�>�(r=<*7�@��='�>V�@�P�}?Q:>�#+����d�D���D���V1ƾg	}��ɓ�/���ͼ��Yý*۴>��>�#��n>�>? �?������>ʕ?Y�?�O�����>����՘=��?���G��F�ξw��=�5=?���/��K�3>�U޾��<��>"tH?�]|��$��q_<�1�>�"���KQ>��r>G/"?۔}��5���>�$ھ�r�?v�i?�#=?��?��<3/�l%��xkb?�q�%���NP��(1��X�aR��4Z�Cp��	7�	��=��ھ)=�%�f>{9>�t;=p|\���?Bb@�:�3?G��+h˾		�B<�>ǳ��v>�](�7Ǚ��x?�	?����>�Z+>$4޾�e�����D�[?�(�󢩾�#�6�F>:�?>�N>rB���~?�:�CiW>�#�=�ߟ��Ӯ�9'=XU!��"�>�*?��=�c">�s�=�YN��3�>�i}>
�Q=~����v>�#8>�:�<lqk�Z ��S��Ծ�(X>�2�>�`J�i�>^}@?uc�?�'>��4>`�?Z� >B��>�����>��O�#�>�c��v�R���9���>s�>��> _=��=�}�G�*lv>G,�>�-��7�>���S�����?`]�>��>!v>9�`?#�?/F >vU=՘���?*o�>	�?�3^�^��EU?���1�?͝Z?d�%?�6>����齽�=�Ϝ>4��O�>q���]h>/ξ��z?��Z�Q?��h�r���U��>��?}�3���l?6I� _8?�P2>DA�>+��D�]?R�{�Z˩<�2�]G��z���b�>��O�O+=�E��ᥑ>�*n�H?���>��?A��?��>9?�B�?s��?S��>�}0�/҈?� ?u\�=��	��Ey?�>e��3Be��䵾��;�}��o��ލ��a�O���!�P��>�"^?j�����۾�Y���eg>��>R�?"I�=V��>>��yP���c־�@��,�$�D�g�傜�+�[�qMB�7��bA��E��6�2����*?��<�wL:��j��k��ߨ$?�*&�V>��?<�)6��q�>M8?e��=\落K���r6>��>r><z1?�z^�峎�5�`�K)F?��e��׾2pY�T�?u�s�<�%?譝�;?fl? �u��?�,������P.�VvE��S�IE���<��-�ϒ��#���]>�_4�>��>������>�̔���>1L������=>z%����m�ݷ��Bp=o��>�_?�W��\?#��>o��==o]�s�J�8s�>���?yRH>�U�>`�D�ҿf��=z��
��B�>��Ҿ�Q��|V��1H��7�??�?*�>ed�䲼m`,��OS?�Ц�)�1>��?å�?+'(?��ľa3<�Ԭ �;L�O�7?�h?�>ɨ> �>>[��>�h����>q��t��e���T3?��?�7Q?�w?T�R?	t��7���ַ���n>�8?"_n?�?9X�=yD�?�w�\�v�92|��΃�k���~��[R�0"/? s�wپ8�����Ӌ�>-C=9���~?ǩ��޺u?���{��>��=' �il(�}D?�ؼ �>������>U��>�>�s�H�h?P,�>��.?��_e/����l�̾�a׾�W?�M �|�Q?��F���`�ʼ_��>��=�����?e�9? �;��>uJ�=�4>�h�<��5?��O��[>�[��X�=�����Ⱦ:B+��V���"��C@>���6>�=����_?y5�>�>�>�k���f����Ľޔ��f���[9��q$����>o���b7��
��QI�>�����P��)�m>��`?���L��+��?��F>�"T?�y�>qk�H��?-ң>Je�>p3l��m5�k��� .�����O?�߻<[3�?o�>/֭=e�Z>�.z>��_����>1pɽ�P����H?&m��v$��������S��`<H?�Y=-��>�;����S��΄>�y@<�\V>���<�a?�.�?���y�?4�?}�?��>"al>�/>���>F��=�hM��)�>j��-����9'��R?��M?�?욄?!�$?�m3?����h��Y��C�*�1❾�5��\S���j��������?�ھJ�|`�>5n<�t[�\O�'����>�)A�û�ɺ����w���a���>���$^��wI�Ҵ?��u=6�>������>�>2Z��.���Xp�?��I>!����Ӿ�?�ϛ>wk�y<�?�7�?Z:�>�U
�+���.&��?M>��?K��=����`>R��>+
�nJ>��>?�{?"��=� �;r��?:���?�qá>I�k=�w�>�Gn<�YJ����� U>�B˾��	�ʚ ���}>qռ<�߄�S%�����=p�\�?��>"?�Qf??��K?�Ķ>7�?���?$6�>�^3?(m�>�^�?`Q?6�>p !?��&���ſ�1�?�ס��pZ�*���ѷ?\Tt�������Qc�>3�<~�B��q ��?��#�4�Q�����ԛ������p-�Z¥>����B�>5N>�=>mQ�){o=羽֩�V-�1W�>������<83>T҅?�ѭ?�B&?�]t�N�>G̲?K:F?3�y��Ж>��վ�u�?ED��#"�n>ƼϾ�}۾Щs>�B�OF�@��F'�D�/��������n?�'�>�X7=G�>[NR�܂�=�t�?'�.?1���@��=!�>�>�?;_���>��?�#�>ۂ�>�?-���s�<>�/�>(���x�]�"�?�j�����V��}�<�>�S�9�[�>��>}X)>��=�Da��2���"?ip���u����w>j�&?mx=�tȿ6�?��?'�G���z����?�W?O�:�W�S?T���[+A>1�<�-"���`�>>[�������Z���&��6Z?���S�\�~:0?˅?���u=,�AA>��_>.��6�>9�?��C� �8	s?��ǽ݌�}�߾�F8�#G/����B/��t��?=>!s��!���y�nH(?��?�l��~� ����>��Խ�����ž� ������!�g �>u��5�)���l�$=*=�}W?L���1�.?��P������f���L?�z4?qP�>�Q�Ù���$�?}}�K0;�R��>�	���F�nUg?�텾}���e>�(�>�,??71�?�VC��dT?U��bQ?�3:�5T?/]�>�J�>D�q�>?��,�*>�3��,>��7���_8�0���ɤb?>�f�<��?}Mƾ:?��>��>5p�>��?�r?2�3?�L>�hq>��0��G>�z<�R���~����<V��?�	�z�='�ξ���<��2>�������=H�#?Q�?�N�?�2?S��>�>��>��(>!�ݽ�[꾷#�T5�EY�>P�F>�"?���}o>d�-?�ċ>����v�?�Lg����>�uN��p�>k4�=⺱��Ƚ��^��t�f?@�?��+�$mJ?��q��N�<� �>y;���澧��=��o>Ԇy?w�>�:?;6��>�'?LZ�?.�`>��<�d<:?�f�>ظ����B�D�ƾ~�U�;�-���R?m⢾q��?W�5�\�M��?��a�'�T��x�>�s�K�+=��l=�'t?���?��=�R�>NX=+��>r����>^�>i��>_�J���ɽ5@��u>���>��'�&P̾�J�����V?4��y]0�*k��_�>�N��&C�����_�?gͺ�TW>�q?����`�3?R��=j߅�<��
h��y��?2	���4�>.O����?�H?� ��6Yz>�d�=2�W����E���*?���>�����@���?d>��=�DD?R��>�Vd�ߥI?��"?Ct?���=��?I�r�8 �=uM��R?�U/���>O�>��v�>yG9�(�>�*���bǼ������ ��!�E��>�P>������>��>��=Fѻ��R?_�����?�d��s?�f���D?����ǩ>��>��?A��� ?v�ƾ}��>�&k>��>�ۤ������ǿ{��Γ><���k"?�tӾ�N?���b]^�c��?�]:���޽E��BZ�<�pg�R�%�l[�;���>�Dؾ흍��4T��p>\��=}n[?vi0?4��>_��>e|�>�v�>���>�?��#�ï_>V�ҿV��?���?�<?[�^?�˄�օ?m�G�����_j�>�?����F;?8�,�c�??��>�2?��?��8?���>^)�?���>�����I�Z<�����M�4?�r��O>�}�?`�h>��?�v1?_RL��$P?�f��)ＫL�����>���=�f2?Q�Ծ��;��G�<b��>�UU�:�H?�g>eJN��&?/P�н==~VJ?�?���?έv��iپS�ľ��+���?�g���<&�]�՛Ͽ��m>��#2?=2����>}V�KB��z�=n�><�0�S��?O0��|�M�&S`��ſ���;O���o�=E�A?Z�
�>P��쭙�Ee)����>��H�Z����E����>�򊾵�>��/��H�?W�?�n(?���>����D�ɾ u[?M��?�=|���,g���v���[b�+���[�>u��>c�?a������?P���=�ξ88>�rc�eX>��b܁<B��y<?q&���T�>A�$��x>?2V�=�#�>����"�>o!\>��>R;�=ˉ?���>�Y�=�ڨ���+=��`?�%�>)�߾w��a��Oi!?K}��%�,?j]�!���Y?�Ց>�7?q 0��I�����%w�?�u��پ�v>�Ҥ>UO!>�X4��l��1�1��_����8�|�����(��<���2?x�������e>��z>��j�ѽB�5?"�L���>��9?��)?c����.����<?�Nn?q:=(J������=�묧>�����5>>U?��ƽ�n9��ŵ��
-?���>���=��k�`�c��>���6�H�H�I>Pyj?��a?�M ?�
�>\��=t�+���ȿM4=�i�?^ɿ}�>���������~?��¿�B���3�?�;��́??�C#�w��6ξ�3z��{�>���>�'�?j�=/�W������ü��9������:��a��`�žL?N��?f�&=_k? �?���>�]h�X��Qr?�?�P<���>w5?��H�ܒ�>��=_dL�P�R���>�۽5E���/>	=�6W��J\>�2�>B,�,�4�YS	�#���;��?�Cx�����\����y?��J��I|>���>���=��b�)��>F��>V���>?��/�Lf@�]gԾbn��?�.����?�"3�6B	?��>?�N�솵��h�?\�O�
i^����?��>�(��?�(�=���8��A�#ʾYr~>�?6�>���Qx��d'���=��������Wн�b?䦢>_YB?�#?>UX==���_*>6@�<4�>�>��¿��>����'��=M����
���;��.����PҾ�>�>y&T>�
l>{�.?�'>"u�>�T�����L�>U�S��(�����<4w��\�Kl{?5��=�U���Z�>C-�
�l�[�>	v>��z��Ƽ��]ȽoPF?:�>?K�T���w��s�ۅ)?�^i>�ȾUX�>O>G���o?�?���vJ�N�\?DwϾ�O½V�2?����NHB>~Z��P��j-`��10�>�۽����1Z�������������2���2�Bdk���8�k�>�I��4��E?>ró���<�le���������ɾˋ���|:?a'��u�P�̿��L�Pq>��>�*��24>���9}?f�ھ�%6�n@$>�>���֊e�O���u*�rk�=��K�����X1��`־����`�[>I֬������qq>�b���3QA���Ӿ�J������>����>��?��?�(=�ſ��b��
a��Z>�7 ��v=������>֓F>�n��d��>h�/������P>�W?��S?�&˻���>'M�=�JJ>�-��F���z>��/�QIb>��S?uL��`?j�>m��?N��>* ?�N����>*�1�;�+� ��`�����)>��D>Ns뽧��<]i�=���>t�u�mڿ=��x�t��?>1<?��>����%��>�X�>r4����;?��I?���>�*��q��>��?I�3?v6�>
>ki���s>cL���ȿ|c�>BU??W�)?P1>�*�?bt<?�N!�C�T�l�l>!���Л>�wD�93L���9�5hZ?�->Jǩ?8�D>pϰ�g�>��>F����l$����X���	����>��k?$�(>�������7~�C}�=�sϾ�J���\�=�*>�!ξ���vn#��{�����������:�lN�5Iy�_;���' >�C���M	�G�;��9JK�][��R��|q������ka2�Мڼ�D��f�>`N�Sƽ�Y#�1sn�O��=�]�>1E<1�u?2k��X�������?Lpk>a)i?T��?3��>ŎT?��?^.�?��S?���?gu�?NmI?��?+�?3X�?��o?��>��_?o<�=1>�S?�1�VR�>/�j>%�I�n���H�>��U�9Y�?w��>!)����?=�ȿ�>q��=Ş��d�݅r>ޔ���^�$��;i�=:��>a���Ⱦ2��> ��<�2�>9eѾ)��?a���l9��{?Zc`��=>�7l?>��K?箁>���g���?��>4��?*�>8$?p~�?ѵ�>"4��+�=�|G�+�B������=?`�>��ʾw��>&ֽȱ(�O�F��-1�IB?�e��?s?ēݽc-<tw�i�!��(:��6?�M�K�ľ��>rJM�v�x�&s�w��ii?������,�?��ۿ��"?�b�>]q?nU���!��Qu=?�t�?RBX�������??����K���=�R��������k>���>=0�>*u-���|<�ܰ= �>�/H>Y��>�2V=(s�J$�>d!�;�}���ۿߝ�b���=?�>��>F	�=Ge��=�`�-�/����?��4?���>9U1�z�>��������m?1F�a��>{+?��>E�ٿ�lʽ9t��R�>�>˾�|ż��>0t~�rF��߫R?�x>?�磾yk���]>JS?��=׫Ǿe�?�k���"�?C�>bC?��߽zH����꾆#"�hp�<,��>�M��V���>g?�k��3�]�
>��>;�7�.�>X6����>�x��4����dI>O��>�>��C?�w�?C��>��?w)?X#��]~f�o}0�� ��{@�>[�!�3��=Щ��+�>��W?�A�<uׁ?�?��"�n�sX>��4�>{B�> �W��Hq>M�?z�:X��>�B�]�>���=�_��A=���B�V��=��־�w�? �ͼ:�M��>5�E�G�&?�M�?�v��j�?>򒾓�>������?7��>铎�r�A>Y�#�-���H��?E���?3��jw=>x��>�)�=���>��[��d`?V��>BZ�>�
R��2�=��>�����g�K��! ?<��>X�)>��l���G?�'$?�	=��ϸ����?%�ν;�ȽS43��&R=2f�b|>C���Ƒ,?�?¾,:����>��E�U�~��z�K^��&������2��u��>w?2A>��ڿa4N?��L��q>m�@����?Qq�?
^�>J�A?{Ҿv�`?�A�>���>��>K?r�<��>0/p���?W��>��#?�(�A}��!����n?�1����5� ܾR4,>ut��w�Z���I������>^���-?���>��,���?Z?��>�$=y��>M>�FξeF��Y�>V��>��Z�0����@���������R���\�� �<��(��o3?�P>4�P��g?�?!I=V��>u�==\�>mu>?��?�5%>�I?�>�RԾG�?bή�L>�9����=���s��>(���0�>#~)�HG>Y���E�����ž� ��X7�8�N��j�
>�a���>�>�?d�L�'���H�?ݸE?%�&>�¾����??0�!?i��>$�=<|�>3bڽI�Ͼǻ"��d�=U�j=ݯ,����ˇv>r�?!};�qb����>�ޔ��N���K�=���0*?\>�r>wM̽P�h>�ݨ�$3Ҿ���?ϕp?��3?b�.?��q�>�>�=A{�e����žq����B�;��prh=1Չ��t>m~���*T�W�T�M]a>�w�>�-{�j>���>ںt>�{���(�>���W����Miݾ6H��*�Ļ��??��>�kO=3�o�S��2�?)�U�;�w���)
>�r��3���`�>� �>�?��Ӿ�ss?�9�>;�>#�����s��>�Ϸ��4影M�>2|?~۷���=��K�]Ή>ȥ=�����S�x�>�	Žw�`���J�Z6����(R���ʾ��������>���>gﹾSa�4����b����eѾ��d?��>9˾��1�c!��E�>yÝ� 睾�;�T�A~F?bHK�V��=vZ����IU��y��̻=�R�$���S(�>�׼=��=?��?`�?>kL?�gI�������;��>T����m=�A?��?z�?�*��u�=��6�8��lE�?sH�>�k����^K���o?ck�R�j?�q?u���tо�#��(K?����5��i�v�?�`����= �>r�?��Q=�S1��!�>�?wYV?�d?��? ->��)?E2J��Eu>���<O`�R�?	Τ�{ ?���>.B����"��*?e�'>
%>Fl�?�ȼ�,I���Ծ{����B?�	��0�?���=�F? Z��+�m>Ǆ�H�ͽ�	���ǾwmK�r��Sە�v�.���>��!>�$��L�D�b?�4���	�Rg���Q�}��~?n׳=@�d>�",>d��>�Y��ҏ��ބ�<������I�a��#	��稾�%R����� �վJ�2����=P��?t*2��Ҿ�� ?Ć�=�s�����%�-�w>c�>�u����ҾԹ�=�Up�{�>�����}�>Y��=+�d�9�S��?�=�j�<��x�4rH���>��*= 3�ʌ>Q�>��>-w�?=�?��>�;���<'������\=��ľѡ���I�uБ>�I���5�b�}>U>�*���=�t2���>����^�<e[�=�Od<V/a�
~.����)�=W����<���ĩ�>޾(b�S��>�0�+aǾ��b��9�>`�z>���?�3 ?���>!������=�vu=];=P^>�=�w˿9���*���L�m� ��%�>��v>�.-��}�/k��*-���0��RJ=�|��Ӝ<�W=E�m�g�C�e����7J>A�^�|�=�&�*Σ��uD�㌾�N"?ځ�>5=-?�ܽ��?���><��>�`�������K?-'�>:4A��]��{w��"fS��4�?V��>�xN?�`���+�����ȫ��mF�,�ᾼ��>֗���ݿƼQ��H�>��}?%kW�Q��U߀>�U$�#d��B�=�5u��N�=��R?��>��>!j��!u����f=�w8�⢅���>&_�>�,��7����珿,��G�Y���n>;�? c�핳���~?ꟑ?�.�����n�j-��S"�B�?:Y�S\�����>B��� ��>�5>*�8���м�[>�WĽ s!�_S����>�tܾ<�n���4��v�>�O��'�x��>�C>�����9�������>����S���˿s ?'1,��m��VYN�Gg�>O��>+��mޱ;)��X	?�v��6?gr�>�':?�"?�8`���?��B?�hu���>"�u>4�*?ҹ���#�<w�>X��?6!>g6^>x,8��">����Ƙ ��Qn��j>�?p:?D	�!ؾ�������D��;U�>�H�=vu�>o�>}i?7�D?�܊?�4�>Q�(?�ݻ;��
f#>]B>�i?���>�0��m�����L?��=����4-���D�>xB-��A?�KS;:<&����J��>I�?�>&?{���$Z;��ܾ�#ʼ�z��2�>�D����bMu=��L?��c�&�b�8����n�>G��J�>=v'��p�aS��QB����?O�V��s1���q+�?��Ⱦtzc��Ά>�{�?
�鼆4ݽI�?�P�?��I>J9�>5(c?��=K��n� ?;����[C�Pp����� ���% � �%)>���f�ྕ@?��?�A@?��.?NϾ� ����>�d?b��>��	?�'�?��#?��p>��+������|�?Xo�=tz�>:���:fO?ăQ���=Z$��龩<4>�^?]����Y��
���ھq�eP���^�>��Z?�g?1y?[�>I6�?)o�?�?��:?�ל?h?K��>��>��?��?b4�JÈ>F;�>&�?K�2���>5[O=�3?GT��t$??>/?gB#�.ҧ��|��n��o8��-��9���ޯ=�S$����e��><�*>�O��5
��fw?W\�>4N��1�n�����?���
�V�T>�]�>	[H���P>��<ЌL?0�>8�y>��p><q����3>�O�����Ӓ��3��>��0>{H���w�l7�S1	�Z��>=@�=��=�ˬ�LU�<!k��R��cվ�@?2�p??{�\#-?���>+�b�
�Z?�f�>D?��u3G>��=��>�(�c�n?��鼏��>�����1�>u�%��ۦ=��=ݸ1?֤<��-?�R�>�~?�>u�=?g�s>��*��n&=;$>��>5K0��Ik�	�.�xu�>[�!>V��L���� ?��}?X٢�^��-�R>�g>���<�>����;z�'>���<�镾.��?���"���q���9>ث��,E�[l�O����>Z����?~��>�Y�>������O?�/�?|�;�*�n�>���>:q2��g��3ܾ���G|��s�(�=8ƾR�'>��<��&�>�2�>ޠ�ct���=ُ�����F���8g>�B\�!�4�'ɾ^�>�����E�G'H>��wM�<�9?ݍs>�Y�Y�*�����\Q�R����i�>�5e���>Z�?�+Ƽ����ʽ��q\?h��>��_b�?q2>�f��U?�@�>�|x�|�=?u�=�.
>IHC?���>ax�?z�v>��)?(OW�>�s��]�>� ?��`��� ?���>�p�=�&o��+�z�׾w\(�����qiվ�8���>`Ⱦ�Ⱦrc?G� �$߯���A?���?��> =�X�>O0�k��Ħ��8>(/���Ǿ�S�=�i?	�1?(7�=I�X��G?�A�=GYP��MԾ���>�D�>��@>��P?b��>�FR=�୾��j���=��>�1K���W?����?���,��ד�: >=�J��(d+?�ߋ��1�?a������~c�>a�,�nP"�=��>lP�>H�����=���k�ݾ�1������jÿ[���?۟>~�~�Ofs���L?H3=�=�>��K�Y�C?d�=T!�>�����~��`�>i�>@u�T)��vi>�D'���B(m��)U?[]x�4��/�~�-��>b���=r�йB><k��J�>g4'>��:����������>��>�ed�o��?ll>�����C=1��>�r���a�'��>��?��x>�gm�����7���?�Ն>�^E��/I�6 J>��4��g��}���19a>7��>��4��9�����<9�t�*��=[^�>�n�J��u��<��O=9B˽b���jL���<=�m�����=�᫽�ϴ=�bQ?��>�Wb>T�>CoR>���<��>�ҋ=�er>�6:=#\M>������W=����XT���`�fY�wzW<'6����.>�߾�Ĭ��J�S��>U��u`�բ��9�>�n�>�M�=~֍>U�>F5K>�ģ�0��JXԾ6��>���=Dk>���J>�	�=-�>W�˾�V �Ow<z����d�����v�򾰏���K��e�>��1>�U9� 󷾆�v<��2>p�)=�Z�FQK=� a<��u����=��_=s+�=/��>�=P)8�({�=�=T�#��9��׾�\��!*>o�ٽ�׽�`�=l�:򥾕��� <�D=w�C�8��=����^��A>��<�F>�9�>�?��>�i�>�E�?T��������/>E�P�p�Y�Ӵ��b�=�Ł�O���7z?��≾�<�Sr�`�[���g!�>�O>Q��>O��>:+��j�6>�/>DFT�����<��*�渟=M�����=��=��=�<�= [S>0�>����	��^��=ox>}�,<�^����=vk>�{���>%f߽�?>�<���������D���oK>��>Z~>��i����=�3_>�v�;Y��=5��=�H>W>S�������f��`�V�jA>1��=�,�;�����=�~�=t����Iμ�S�;t��=�BԽ�~���?gIF>mw�>���ƪY>`<D��A>������>��z>�">�R�L[O�����*�R��릾�c��i�1���|��	��<�I>3��=��#>K�{��ҡ>2��=��>oc���3�=L�>�N�=Y������>*��>R�>E��>H-�>*$���$"������{}>^ƽ�e|��O��ú>��q<�=&��������<r#X>��>/��>;�U��4>�A�<�v?� ��L'>��> �>Q�>�/�m.�>�?B�
>O4�>'�$>{b�>�E��v�@=�#��Gi�>�
��ߧ���|Ͼ���>N]�z}-=���<坶>e����0?��"?܈>�-�Y*u>��p=�!3>�5��;>�Ȱ��.�>���@mu=�2���9=��<�'w�ά���ľf�<��V>ܗx��|5�
m>	ϔ>=�s=������`���:>��T=�.2?-�G� "�>�<����>�Ѥ=��>BϾSB'�ɷ�=�g�����~��=rf��9SM�}ߡ��F𾖀c<�F?�<�=��>�W��=�O>z��I�~��>���xH1>�9�����M����XQ����=�<-=�D�>�9��z$�4��0֩>��,��1��|���k=�HL=>5����g=3o�>����έ,>�-C>;��>�����v<�ǃ���t>݈پ��=�=.�:�����;k�9-��v��<u�%��&!98��p�=&���;�*ӽ��=1�8��������0��=�Y=q�=�W��Z>;�νf��(Ť����=�r�=,9d��_=�ާ�	���?�=�ݗ��z�=�v�>y?l��>��>W�P���޾Cٟ���=��;�{�<�\�=���<�~�L׎=���<��>��z>��>��>�\�>C��ຼ�^����=e�=	NJ<�P���d�<�>�d��u0�j�
>� �>��|>[�>��9>��?/�>��>x]O�k�=��ν��������.>3@�������=N�ԝ��P`��т������D������'��=?E�B��y��Ѿ^�?P'�=e�	>��ӾV9=>-R���y�<�n����=���>ܩ�;}�>���9�>�X���S�;��I>�A��̫>@�Ͻ�k���7�������S��O6>S��>��>��J'��М�=��,�� >�<*>h$=B��=���v�e��oξ�߅�������=�����V���<w�}>6R������,�<��>遽�W7u���0�u�>���S��=����k;%>�ZK�`a9�Q=�>*3���yA�M>�e�2�þs����>e>���=H���=۾q�K=�*W�ߚM>S�3����=�SA��f>�W�=b3�T�p=5rg>���>h�?W��>���>��@>�?!.>�3>��=	�>�R�����=�Vk>�ͫ��<>i ��>@����j�[�Z]���^>�̀>�s>��=�Y�=[1?��=�>�=�X�=\_�>d�ʽF8=�fA>��t�K�R>��>�bh�ޒ
��лU3v���`>���\%�>��-<�ֶ<�P�>���<�">�E�>�J�>��>@�>K5�)K�Tc�ʆ�6m�>��X�JIS�7޾Qb?c�����R�-v�=h��~柼&��!����Pu= `>�ݝ>��Ǿ�{�m4��M!>��:#��fW��h@�=��l����#~��<�>�D�e��=|�>�D�<!�þ9d=���<&	>�����Q7>~'u>�_t=������G�x�O�J1��'�)?��c?Q��>kk�>[Z�>A��>�a����=�/�>_���l�>!�>uV��:��X��m�=��0I?Q�=���>zI��$A?���<8�y>+ _�w�p>��y>�n>S�:����굽�Ǥ�d�@��?,��>.��>�}=u��?
�>l�X>b}R>֬6?��>;��>�ё>w�>Z�>�'�>	y>G�M�-	��?\DW�v(S���'>
&=0��=�ԩ�� �>����>��̾U���Q̼���=d���ґM������4�����]�={ͽf�[�Yj�<1|�=�� >1�<�[�1��������g�E>�P>M�;�&���;�=͘?��7=Zù=�Y<x�^>�n���t����>$*��nX�=�yG�i|��Rg�xw�0�p�&�9��
����<O9��vX���l�=����]��R>��>x�=�Z+>�ؚ>���;��=������>�9�=���>�s��;�=J�
>慂>�䈾��?��=޴��M��tC<�)�[��}��k���1�<d:��A=����ڙY�B>H�=��z���n�Z>��=;�5t��׾S�>���<@�Z��&Ӿ�O`>���>̗=��R��>��>/%�����6D�=}���`f~=��U�������=�)�>�����;����=�Rf�(������ �����=�o޽�#�=��/�,>s4/��h%����>H=�=��-�t�7=&S{=�h��޾�ƀ>�`F���;>�0۾�wI�n�S�	AV�Do����m�0H
?�n�=��߾�����=}���v�����=�ޛ��=b	��}y�B��������۽N.�Q�꽊�Z�W{�>���='�=h�����M=�Ia�[�f>��>d��>G~5>��>�;�w�Ͻ�Ps���=�Խ�Y�=�d=��>��5j�J��)=S�]>��>-�?w�>�.�>δp?^� >�c�>��`�=��>�^�=<��=�)���=G���h>��}=����A����iy��i�������u��t�������^�>�9v�^A�<�,E���.>VO�=CM>�����I=���A�<�ν��������9�1���>Y"켓=u��m�=l���d�=���>�B�>zH�>���>�'�>`��>p�9>W�>�3y>�pa��T���o���9>���p����x�8�f>-�eM������w��>DM��4�_�xY��N�x=:H��W�~��OѾ���J�L>Ҷ��.��{��r�k�/��8�b������<�8�'�ŝ��GՀ>Y砺�ޟ<��P=��>�b9><�T>�f�g����7�=5oA� ����3�T��K��B�;$�<�C�>��g���;�S�a�=P7�=�����`<�1���)�<T��>�{?�T�>�?�ږ>3�������=+�>w@ӽҢ|� �]=��>/�������=�Y�>4�%�8�ѾJn����X?�����ѣ<�=���?K��DY��5j��P�>�T1��q>��$E(>�}�f�1?������*�[S?LԾ�{N>�D��w�>�q�S����>60���nY>4l־]G?�z?F�=�_�>$	�>�Ll>u�?�9�?��%?�����J>�1�>D��>��WfL>��>]ɽ!��"G�t�>��;>=����ZF�3���!
�7l?�$J�c,�>��>?�_�>ih��?�Z����>_n�>�ܽkc�����>�?�=���?$�g�Gm?���>���>H���h��>`)�=o�¿����ݱ��.��]ڈ�c�X>S5?n����H��.�)����7�a>����q�j?^cK��t>V}?v�"=��>>m?������uk��Ѥ�����|P���V���x�e">e���2��>���>.+G�+2�?��z<����Ѻ�"�4?�Y?[[�=��������J?>��?9�?%��?ݭ�?�/�����=����*Ӽ���M�H�O+�K�J>�+\�	���\����=�����?��|ÿ52�36P?���>��PC?����Ĥ�A>>���>bV>�������u���D%��t�Ҿs���
���?���$Fm?���[8ȾmN�?�м��N
?��þO:?="����,]?{5��:hH?n|�<'�5>�!�L>�N?�z��x`>lL�SE�>Q���8ط>�d?h�:?M)?myþߗ�>�/?:9���i���W�� �C�?̖�?�N�=�I��bT?���=6S?~�d??�`��U?��S?֓��cW�>���?l�g���>��?Ϫ?�K>V@��9�0����">]K����?��~�v����(�Cr���ʿaB#?��Y<��D?Y�����:j>˦P?�4��P�9�d��;�A���a� ��=,�S�E��> *P��wl��v�=��8>о�?I�;��3��c�>�8��n>J�m���z6<�c�>��P���j?|��>�����e��̌�?�����i<ߥ����?}C!��fN?r>Ž��>?�77?O4�>BT�>����IͿIӽ>�>5i
?�yܾ�V�����=�O	>J���gu��?b��B�g?W�����>?8��	O�?�
��V���?��j:�?���?��ξ�`���5U=�Y>oھ�%v�7uO����ɝԿ�)�o^���DZ>F��$ſڦ���T����>�^������@z����䶰�q�>���?��	?4u��c�%=���>�P�>�.�?X=�<?�[��P���g��y>�<<�:���w>��=q��>�;��?$�����?��=�+�o<�>u�?�>?e
?S"u�53=����r��2h���?�W��E�z�=ַ��ω>	���.[þ�_�����^)�R	> A��(�>�lU?4v�?�?�P�?���m�@���!���>\U�=�q��.����G�������>'���'n�f���U�=q������>F�f�� �:ДJ�p�>EfW� Q���{�%=F>�j�>�s
�C�G?�'�>����"Q?/���K��>���>�q?����؎�C�]>�CD�ՠ�>����V=�!>�MA�VXP�L���T=�I>�4=�p4�"un>���;�o�>UQ��`��s��e��(J�-B?d��>|;<�i����>�1���u�Y$��P�ɾ�,��.�X>+@���/]���W�y?�]g?�m�? ��?)Ɏ>��?�o�?Uf`?�6��O'�?������=�9k?��D?ܞ:;�p����>�s�?�o?��>G������b�ξ��D=%?�W?}�r'e>�0��m�������Y?��Ѿɛ:���n?*?��p?�Z�>P�{��@"��' ?�*?�hc�:��=C�>���?R!�?�ص��:�>ׅ����\���͚N���?J$\�ص5>E�J���\Y�i�M?��?j�?(��?[}����?�l�?WX?t�>1�>$P�=��g���оs���`x������̮��pv��!���a�D��>��=T�����;��*>�F>j௾[�_�b5��س7��ur�R��K<ɾk2;VC��2@��q�=hǣ>=Ω�dO��<?J+�?�O�=�Z�����_.?�+��h�����Ֆ��i�=��>��侖Gv���Y����Zj��L?���?g?��?��<>RKؾ8|}�U�q��.�?\	g?2��Q���Y��Oɦ��<��n��~g�T@?�24�� �U4?[I߽و%?�N=��?�Ψ��k�X�?e��>#P�?.�W�g��>ȁ���v?q��]���da?3G?�¹>�󌿢
��s>��?Q����D?�?�>��>x<�Jj>tO��d�o>֩,>��g�!��҈����W>�:]>
Q���8>_�5���ý=>�������X����:?���`��?u5W?�?�O������?��=?>@���zs�?!i߿�M?��$?��m?y�Q> O�?�#�>�#?���v�>Nu&��*%?}�����? A�?��˾)��ί)?��c���>�e>[9���n>��]?h?�[;K�J����>�!�?��?°K>x�>����Έ�x�h�¾���=����E�?P0�z��>���>���?):7���?Y\�i�?{C������xd�(O">qz��Q�>h�X?��?k<l?��m?���>�i�>EN?n��?��l?"��?r�>�1�?z��?3�\?W�?G���?n�<��V?���}"?UA-�z�>�("�e�p?���>�*h��I��J?�s�������@���~=">�f�l�S�.?�>����齄>Q�L?���=p��>�*ʾ\���e �f྾�k���)�?�u�e;�]�>�(
��>�m?R��>o-�T�8?�2^?�N<���?y'��0?�.��6=�����pR�k�=sZ?*�������������>ZGI=�E?R�W?{A?`�?/`!�7�;��2>F�後c��R���w�>�/1����>�W�� �>Ѯ۾`����-�u��=T�ľ�(�̲����>��;=���>��3>�XR���>�˅����=�By?���>��?iY��.�?���g8��Ǆb?����G��
ח�73�>K-���QL>̝����?������>�B�rxm?�.p?&8�QJ�>x_3�E�K?�g ��u���K?-�K�m�A?�X���>2]�7��	,�>���c�>��_�d��PF�?,����s?��0?U2d�U�п��>^�U?�T'?��s?����
�<}B�>�Ӽ��>.�P���?��~����gD�>� p��6��߸�> ;�>3��#m�?}�a�ǩ
><����A�M`(�e}�?1��6B�����>�������`p�==ξ���>Ǐ�?���� >�:ǽ���>�H��4��=��=�Y��	�`�J�:�>�S��G��;�����>��EٸpsK>Tt���H?o(?�b��C̾5��=Oii?����f�<�f�>��? �Vu�?�����?��I�	��s������W�?2�� �=36?>j]��">���?������_��c?;7�?��?�p�>�W%?)](?�i�C{������'�-����)�z��>~M�>6��><S>gMN���-�?��>�dz?6�?���?��	?�$��L���'o�%gA��'�`������=
;��W?��J?�	8��\�]���G� ��8ّ�i9�> B���9?�4<6<>z=*�S�ܾ�f6����lȾ�t{�_�j=��?Ed���]�<��)�w �>3q<?�j[?}�ԾkI?��?C��?�uV>�&H?`�<?]b�>'Ρ?�~�>���>5,���f<�Z�=b>D�">S�>�>���>�.?»ؼDď>�!,?+�?��c���#=�u?��>Kj%>���>�E>�I��>�-�)�-��Z�?t�=����?%8 �k�=��ʳ>�q>`ԓ����>��Z?�	/���X=����d�=������?�7��O;[>[�d>B<?��Ŀҙ���1?�?k$Q��'�>x3
?�3�=��ʻ=��=�F�=r��;lt�<��;h��~2�r�>J��ߎ�;�>���Ľ~�T����a�>��>�@$>�>X��=�\�>�j4�?1�ܳ=�<���=i���
N�����[��Y�S&�<7~��6�j�=��p=��?�̥���j4>`.ռ]�x�#%�)�;>0΅>�Bd>��[>I*L>,qh�"Ww��wx<5;t�ϝA��=
��<�-N�^L�<OB�=��	>��C��Ǯ�r����$�>]�$1���n�������������B��=fM�=�u��2�=�5>3�2>�3��p<��7<�k��>�ǵ<��=�`;>ډ�=8���Iyݽ|ai�G�S=�>��^��*�<9��=,�<�F�@=|��=S4�+���Gd=����}�߽�0����<юo=��ǽ�:��ڕ�bz�S��=�DE>.�=�	>M(�ǋ½�#ٽ����
<��Y�<�.�w޽sC�݋=�"Hs����<h�g��0��m���@���f>�'>��>4v>�C
>���+ꍻ��V�:�=ܽ �3���p�)�%��<kL{<̳�=�c<i��=�|w;��>��=�k<�ʀ�m0�=%����D��u�����;z=�����ս�X޽	ӓ���%�И�7�J�ؖ��WF�'�F=��>&t��OE�ؒ"�e��<(O��x�Ž�,:�޽r���BD���(�[��a���G�-ּ�Ϳ���o�_�A=Τq=�50>�+�=�В�_�ɒ����k=��<8�:>�3��Gc�	M	>��=?u��W�>�Wa=�Q>u����m��e�����	t��x1<5#C=?�}���@�A5�=����%���ҽ��=���=OPg��`��b��6�=�����=}�W>#x�=Y�@>��
>J{�<�l��Z��P�9<1�B���:��3�<�e�}����ŽDi=�v��_z���>�`���d���н���=pM�=S�M<�ђ;���>|��=sг=x�>�#B>+�)>��O=���=;3>�!>��=3��=8"�=�̽r��c�-�)J>�v<n�=>�>�:��e>�>S��j>I��=cx=\������=_	2>�'!<��Ľp��<����A�>��}�Xk/�:U����<�L��c.���ѽ������Pܠ�Ǔ+�}[�<��j�)�&=�Q�=���):���5=z�4>����=>.gc>�A�L}>�0�=����O��E�Uy;�V�<T X�!I��Ixӽ��i���(��<���Ji�����u��<�m�Z�=Rt=?� =���gMI=u5\=��=W���>����Lg�<Ȑ>\��NO����=Au��� 
�*�+��=�<לĽ]��B�]� >�=�>݇���6>)��=��>/�	>�&>���<�=p�����M/�>L�Ǳ���_�=�Ž�c=���4�n���&>nS�=\!�=d��=6�m=��q��;�hQ�jɜ���6�a��� �=ɓ�=ٴ�=d;��>�g�y@���ż�ٽHg�;�^�<;�U=��<=o��;�)
����d�at>���>�2>H�:> e���	�}p">�B<K���K��`�=�#>:g2<�d]��tĽ𰮼?�>՗g>�(S>�b>��>�=���d=tKH=��$�gxܼ��g���6�F(���%��=߷�=!>r�->�C>�C�=&�"��a�j0�=m�;qϭ>��y��u��ry�=a������=��^�A��$5��D��G���(����'��?��o 1�ɼ�
y=r3�ʲ	�2�ƽ�_N=Ե���H>� -���*�;�R�ԅ>=�sd=��)>�l3>.N��1N�>�@載I��*�L=�q=��>�O�=����ټ�	�rӼ��^_;�3=L�½X̼nq#���%��K=��j���K���n+�X�}=E���G�I��s��"a�#��� �o>^��<�(?�I4w=��8>�_��s⚽*#�+>�ʁ�b�c�T�<9�L>q1�=�ǵ=P'>�ڜ=�6��T�VN�B�=*S �T]&�7n�t�_=>�"�v���}��w�>
溼}�R��?�<���)��=U�ht>nK~�:X�$ۮ=7<�=�}ͽr��a�(��=r>b�i>H� >Һ>���=���=�%=�>b�f=�,>�Ѽ<�����#1=�I�=�ȓ=�ߵ=v*Y�R!g�HXɽG�+����i⼘�)����N�;�������
��=3, =��;�H�.=9�o<��܇;fz=��b�,���+�=<>�E�{�ڽ��=H����x�=um=����<GWؽ��=��>�%>k.>~x%>WZ����;��G��9��*Z��{�����b���P�i�y���1a��ٯ_=��Z��H�?a��>>��:>L�y>�C�#���Pu=z��=�~�Ј���ҹ��[)>C�����<�a+=$�>�3� '=��=�+>�\B��>�=%�=��>6er�Ą�=��=vԀ=9�8�p�`�4�������B>[X�=E��=PK>�H�=�A�>���ڙ�z2�=}K]=j6>iV>=��k�f���$<�N��<)����+
>�Z����=/�">d�<�PN��.���>���=�v ��(���j���2�!�F���>h)>z=>!�=v>7jr>�g�>���=l-�>#j>�e>n>T�?�}@>�\>��$>[,@�J&��&�2��=ĕb�5R��a�9=�;	>�R��!�9��=�Zf=�s��! ��c��.6���>���׽�$�����ۢ����=���<w�<[����=�&>�/��	�^�ȼUꤼ5]�c6���*�����Y��=��=y�\�v$=��>�#�<��=~���>Q�e=�
�=g�c=��D=L,>Z���u��v�$=s�l����=���MO�=�~e��� ��]'��"W>t�[>���<K��=���=t)��̨=�E�������>,�R=���aJ��\�=�h�>�ѽ���<���#��,�H���-�<j��E�׽�Ǽ�s>>*L�=�Jw�<�7=��=�Z1>��񻵂Q��ƫ=�~�=��$�m/,�g������� =(3�b�r�K)�=��#>�t1�p#A=���=��=�����ޝ������:���{ >�n)>���=�%=c�=BD�tt�=�(ݼM�½�є�rM��t=�m����O�=���� ����:T�׽Z��=-��@�P��E>^��=��0����<꡺��>�(�0T��N���4;)k6���������U�-E�����~�b=G��<���Ҍ�4=�'�׶����r����}.�>g�=�Q�C�N�Ă��|`n�Z�,����_�=�=|�=52)>.�>>��p>��>]>�	�� ���Z�8��<oмL�)�n��=��?>W��Ͷv�N�=s`>�ی>�\w>�Y>?�>�W\��|�=1�">y��F;>j�=�8<�[i�敬�zQ�=��+>��]�;����μ��~�̘>����Df���N=�f��� >��=��=-�;Ӽ9>�F�>1G>�A��(��<*½�4<�<��&X=\<[qӽd`����ʽ|�`<���=� ��R�����m��v�M>G!+>��1>D4c<U_>��4>,��=��=R=�W��u�:��A�8��s���a�ѫ��Ȩ���-�Is�<^�N��U;95=�
=��p�� >��S<+Lc���}��8i�
m�;R�;h�D�{k0��ͽYPR�O,����}���=�+�t�L�j��=	��<��=EyͼU�=��=��=<���34=b�ݼ��1�i�b�4���]@��[��[��q8�<�0Ͻg��=�d�M�Z=�'c>P�>�j����b<�>��f5>��t>q1�>�:>mַ>P��=�K�=�E>[��=�a�=5����X�l7	=�=x���sV��2>)����e!���ǅL�Vm=�˽d�k��a�����=���=z˽̈���>��w��%>���fjݿQܾ�������NZ��vϿ���=(��>�]�=�2?���8��{ ���Y��db���>�	�?T��=�8=Y
1��Gg�G��<�{�>T�>��?cP">u�(�A!�>8���.N�>N���8��]����>�x�=�=tK��ͽ����僧��w0=���>�?V >�nQ?'bt�L!@=��?��w?�j�uE���1�>D�>|����=�
�� X\?D؇��l�Vl��-==�����,,t��@�^ƿ3���e"�^@հ?�sྒྷ���k?���<\�������cu<פ�>sq�>hF=L���/�>�)?����N1����*��(~>V0a>5�=�n1����h-��fdξ(`���%>*�>\=<:"��~}��'�<Z4h���Ӿ#5�>��� �R�>G`?���?�5g?K^�?�O�?M ���!���v���?�-g���:l����	?/�þ�ƣ>���=�V�G�9�Z�
�x���r˨��S?�!�F�=�W�>���f'���0?9��'���J>[e�>ԓC>�����|��?@?�Jſ��0\�=wo	���=6 ����?X<�>8M"?s�2?��@�r9U>Ǧ��&�����P�B?�m�> ��[ ?߆	�*��?�P+�7=.��|�=�*R� �?D�3��*�H�u�� �>5>�4��A���JU���s��׾]��?�r?�9�6D�0TY��뛾P�L�A�-��{ʾn�о�2�>$����������B6T��Ӷ=��ݽ�>�vB>��>ٜ>Nf?bK=j�K�Oq��D�ڹ�<xȽ��=o��ru��hpd���?��
?X[�> X�h�7��E>��>�>'}?��>�b�>5���t��<h���aɾ�?Y�(>W�)���=e�����>���>읿zx>�J��pr>�RW?~3߾�������?�����?"�V���B��f��iY�>�4��{;˾�#>U�?��C?���=��:?=Y?̋�?Lx�>I�=C2?����>�������?��>C[>�1�Q�=X!y��&�����>j�}>�ܬ��'U?ԑQ?>^�<�킾�N+?�"�>e?�eJ�q�@?t�̽���=���Y�y��R���po�K쨿e������_+D�m\;?��>����x��!=�>��I?e!�x�ϽM���d�>6�>� ?��Y=+��>���0e>m�\����� 
=������X���ા���뉞�*�׼l�j�o>FuG?�L�?�dA�t���M�?�=�I�?��y�������?B�L��󀽵s��|�W?�;S>()1�2�>����U?)�?'����+��/>>r���B��f��[@/>	� �<]�h�'��>?^K?'�?��I?	��?����с>Ռ�>��? �j>�r?�����y�>�'�Tyľ�-+>o��>5Ҿ�{Q�cN��H=��� ��=���͢6� {�/�-��Xm�]�>���>|��>	���/6�dt��vv�G�@?lBa?[��>Z:�?שS�T�)>3v�>"Ķ�y�A�j9�=� ?�N>�O�?��0�������Y(?v�>K���C�??�^�=NS'>��c�-?�?��"?8�1<�m"?6�>��!?�k>%�|>��=��ս6���X��p-����Aw>)��T�#D���h>*E,?��>P�>䋐>w+�?�"Z?'��"�<��_��d�����>7yh��G{>3FԾP�>iS����=���7��p�=��+����|k��}�=�.?s���f����d>0�
?�ɿoN ����X�Ž|3C>%����*ᾃ�L>�� ?��>=�>7މ=o���v?lS��Z+>�j�=⯑=NX����F�U�LF�sGﾰ,J>��?�,��+E��c���@��z_>ТA�Hxw�*Z�r>��ѽ�K����j��_�����=XV�"�l=�ƌ�{�="0-=��>��a�@.־+?>��P�y숾��I�>V����x=4�?>
*�>��ܽ� ?��о��|>䓢�j!���P��C>$�^��ɟ;����}J�>�Ԍ=�Z��Z�>�R��#�?)%S?L���=�?-�E���J�1�¾c���w���l">W��o��=p��>�kn>����>g7��$#�)�F=�M�>��M�R}�?�G��$��į�/�Ծ�4�Y���#E��0���/����?E��>V�>xɌ>�>agO?����Bٽ��V�y��?Ӿv�?����Ϗ2?���>�\��،�� ???�T?m��w�>��Z�
�e<�����T�>1������I��>���>�a?U>�P¿א�	j�)�a�(_<�H�9<a���@?�����>l��=�U�=	@��^G	�������ȿ�2��;'��4�?
;�> �&��������><��W�׾.1->5@5>�>ˁ$���?F?S>nX�?��8?��ŭ��!7�X¾r?���>>"�?��;�P_?���H>�1����of>DvT?��dRS?��>��n?��?�Ҙ>>�;?ծ�>�#���sP�|[]����P3���9�>C�ξO*��H�t�ȿs?`���A>��-=�d?�$�����.�=�����r>�H>)�(?=v?k�]?�=��?�]8?>�;?�H?�?��y>�?��~?�v?��u?��?�,3?�Mn�$��>Ήa?b�=Cu߾fR�>��G�>�?�Y��>R/��k�m?�\�5�f�OZ��'?�7�4e���޾r�,�4Y�:��>X	�>)��l����>�>�[ƽjی�;�;���>�k��o\�?lKM?�A�1�=�����Y?c@��IO>��;�8�*�SE?9�о�Z�>��>�F���t�L�>��sk?���G�=�v���G��n����\g@�?�>ψ?M')?�bv?4�U?x��>���?J&�>���F3Ͻg(��?���=�A?<����?�΂��> m��|p>A�>�I�>�D?�,�=�ZG>�v�b�?w��5y�>�[��	:��{k�=_\���������>��>�U
?c#+>φ��B��?�#?ѭ�>񕯿��?<57?��*?��_�=�<>�
�,nf���1�����ۄ<�
���ӿ��ľ̘k=��׾aᦾ>���n�?���>`�>V�-?C������>^���d�{P��4b>�\><�0?k*�?����|j��!�>1��6r1?ǣ'�\_"�X����?e52�LK�Xl���;���0~�ܕ?nY���[&?Q�i
�����>�5	��@�>�Od>|ɋ?,�<7�9�=������@�>�?g���˽e~E�GA�,�\�b�!?���=&s>��W=MD�^l)?�'%?�6��c�#?�U(��q�?�ذ>�y�>D3?V�>���N�)?u�>��<ϲĽN<,>�F��n�=rP-??=�=8��>Jk�>Ti>|����>;w�?�+;> ��=�d2���=?`˽F�<�����G��B��>�辘�=�ju�?��4?�]>H]�?I�y?��=m�>�?ZC"?e�
>�&�>W���Y~?U?h)4�;m��Cu;K�_=::;�Ȍ<u�Q=�����l:��:�����
?��?��A?�8p?���?�x�>ác?�O|>��,?��!?n���*~���E�)>�,�>d�n�ES����>�l?c��>I?���<?�,v��[y>b˵�1F���6��+kܾ�8��cN[�����ܽ>2Cﾭ�;?���>0㨽ζ?����a>�K���EؾBb�>�T-?���>�H���Ɏ>=��>+z?K��P��<��_�r%�>�`j�f���>ϰ?� �Ty��A�>� �>}U�>dΆ�r�V:�>@띿������=�'[���3�un?�k�>�t�>���=k.?�2m���r=%�>k�I?M]=-�
�,�o?��>�Ĵ>L0?[΂�K��>�;��.i(�
�/�S�?�tվ��:��a�霺>�cG�A�>��t�yq>ߍ�>a:ͽ�K���K"�T�����> 0�?��#?L�����>�����?MqP�������=��&?���=��$���.>�@I?�u��)�r=�?��^?��	?�߾|�+#�GQ>=+">?��P?���>���g��(RF�t�T��A?��4<y������q?K�"�����T��W�������D:�e�H>k�>�>$�?5̗?��f?ŧ'?v1{���?x�%>	U�k6O���ﾎn>��m���<����1?��p5��~d?A�J>��)?�)��p���1ؽ��4?���T�Y�Am���uG?�qW?FD?�ľ�T���,H?7����4���?��?��y?�� [i���??��3?�:���1�=�y�>@���~w>�Z=W�A?��?L�����>�6辟AO?:��>�2?ܒ���>=J�=Y^��<�&?ܝ>=;�>P6?E!?�m�=�{5?���?*��?��A>��>�X��?�z?��S>`,=>Y���?�1�=�NL�lʨ�Eh?c�g>�+N;��L��f�� �=>�>º�t� ?�5�>�ё<�s��G�Q?�y?������V?ޟu�����^�=��?��@?��>"E�1��[.B�A��>�f��Z�;>(.���I ?���=J��l��=�F�?�o���\�6?Ui¿p��?J>ҋ�[�q?�^:>>�=6����>u����<@ d>:�J��]�>���ك?Y.��񆿀使�b��m$�X��?�dQ�N$"?�	?�$P���.�t3�!V���,�?e�?N%�?SN�O��=[!�9?��<�ܾ�c�=�����2��sJ�⁪>q�	>��\?@l�>��Y<�����Vӿe�D�e�Z�fL#>-i�?�>)�>5>�P$�ɖ�>*�V��ý�s#>�T�@���S?������n� ��,�>(3�ب>+H��)8�<���=∼,Ó�)@��i�>ӂ���|6>Z���:�;�.�/��Kr=M��
A��
�p�>�b�>P{�<��>&C׽���T�׾���=��k?,2�=�'{?��+���\=��>i��>�oϿK�o>7�"=�ɿ� >���>nș��d�?�c?�|r?Fᚾbv�?"d�>�j?\UM��ڻ?�*Q��������?���Tfk�9S����=�A������m�G}���������=R7Z�p�6��y?=Ɐ?;d��	ľ�?p>��?D��L�W�Lt�?��?vy�>�����_>�
����>�(�>������=�P%>��+?2��8G�C��3��>�\>�u����N?I�r?0�)?�������<C�T>ʠ�>[�Ⱦ����!5��������'�·��w��<� .�$t ����>�4q=�*v��-�� S?
ݓ>���>6m?��>��>���=)���?#�½�?�*>�/J�һZ�,�=���z:8�xU�>�N���n�>S���ѓ��d�<�М���z?v��?2�>�!<z�[�E���'�<�^?�V>H�������r+>�T���W�4�W=�5ؽ�N�t2������Q�U�p�=v>/[?S��=����5��w��S?��?��B?���>/-P�2�o�6�7<�C�M�žwE�=}vp�Sɳ��f�>��i�Ȗ�豓�k��?�ޭ?ӻ>?;Uk?L�>��1��y?��?�?�:���D�Lb��<�&���4�R,>�7];O5��g�>�k?���?4y�>(|=���[��m��Cm{�0z�>�H?���3i�?���+��3�y=�Y6=��I>$3K�cͅ>A��?x��H��<�E���Ɏ�����?g�J����= \y>�e��p�?�6%?V��>�鯿ߠ	�S��>Ѻ=q	?��Z>�#�>ǻ�P�:d���&*�=��M?\�[�ͽ�5+=�@�ĐY���=�u�>ὗ�FZc?.�%�np?�ѓ�Y��>�e��?�m�?�?O?9�U��o�_	�c9?��;{�龳y?�+j?��k?�Ŗ����Jl?'�G?�ľ���>�ɶ>_�?�~�>���>��M?�:)?���>o�?�>���>I��Vd��+�>w�i?"w�>aË?O��>(�k?��t?H�?��`��g�?a�X��˾����)̾����g�>"/��]��>�ƈ��y�?T|�=	>��?��>9d$?6+?�B=���>���?�2��OO�����̆�>�M���ؽJ���EL�� Q�b��Asr��ȶ��bl����>e��� �>�F�;u�T��;���]�>`.�
����%�8�Ϳ�s���o
=Ӏ��(��>�-�=t	?����'�$�)�=���'�������=��������
��>૑>!�?�إ?WTC�h1����>�5�?ӰS�ԟ�>�VE=ԵV�[nu?���?X�!��A�����>���??0?tQV�=`�ƅ�=Rx>v��>������F����?��:�����>�s�<x?�0?�UQ����;ß�=hw%=���>i�6�媾���>=����A?&���j?㥀�J�?Pk�>��� =d�z
�F�=�]��em�}�H>u"0>M��?.�f?�8��#�����>�4��!>�`.=�`X�x&�2_����-�H��=c�> m>�i>>�I��.� ?�R����=�=(�r?wE�>��	�x�Ӽ�듿�aU?�$����B�����%5�����o^Y>k%�=���
�o����B���X�=F�;>[����e�<���=�Ѿ�������Ԛ�?�OZ?ƾ�y��d�I?O�>l�S>�j+�?o9�VP�>��}�|>�F>+��>|�ּO�?�?x"?g޼�|*?B;�?a�%?�*���d	?��T?=�3?�D\?s	?�]�?Q�?3[��{��W@�X->�g�徉OE?��7?�H?�=q �>������>C7�=`p��#]f>���n�f�/��Ե�=�T̽3�T��wS��u�>�  �Y�>;߾��^���>dFN?)�[=��M?c.E?D��>(��?�H-�' ����Ŭ���>����0�?�}�*wZ����ΰ���?���m>Y�پII�T(k�-!��v��
���e��Ͼ[1������վd������<e��3����8����(�>=\q?C�d�d$����œ8?��j?�h���9��뫾&��>��ܾ9 ��������?ͮ�2i��R�6�A�?O+�mG?��~����>��$��pG��۾M3?2���-J?ζ��E��>�/��v�>̖�>���� ����wRp?�ƾ.%U���¾�v����5= o�ef���=�+���j�X���u?_��>ng��0>	���MG4?���T��?fiu�I�?�`4?�&7���ǁ�����a���j�W�'>�R���'���x�?�?׷׽r)�O��>|a%>��J��\�>7Hs?�"�>�R�\ྡ7�?G�?�����T;?񸿉�4�T7?c��j���A��>��i� aｫ֪?��8>����?�+�>6??��<�?c�R?_���b�=�N��)#0�\p�?�{F>���LpL��*?�wL�=�;�܈�Z[�����?׾ef��+ž�39?[I۾��ܾ�'Y>��)?|qݽ(���~���>�="?B*n���m�����/��὿]���ʽ�o)�G��>��>���2�a?�P ?UӁ?�*?�K?�Nw?g8l?���?��&?��-�/�ľ�ޙ=d�?�ٕ=��>~sj���i���+�2��*1�:w>��!=�Ѱ>��>�ø�dx�>�1�=r+>~O���z�?��?ޫ=0?�����5���/�x�b��ha�"g���&?��q�?�l��Ǽ��Ͼ����r��e����s�:�`>�"���<�>r�+>)"?�i��w�=�bž��8?k��5��?���P�?��-�,*g��+�=�녽�u�>'eᾏ�v?�?�1��8�
�#?�	-?_2L��q۾ ��>J0��(7�>椉��iq?M���0�����%E?���������>�V�`�>f���P���e>"��>�-8>�����`?������,?A��+�?[�	?��=�ԭ<�P�N�ҦR���:?�wۿ�����>��ag�>�w����=��P�\[�?� =v�&������
@�m�?v�q�	�@�?��!?�18��b����>���>��V�ڭ�=������?5{">1<?�G���W5� �=R%�?a�3pq��s�>:�><�X��X?ߚ?��>�p^?(xX>�����{�N����˽T+U�QLƾOV������f>H�Ӿ���>R�>�Q}�n]���CB���j��ho�DPg�>錄��)@��?�k�>~����>G�n?�i6�a+���
@dd���?��5����?�����?'m��˞ӿ�l>@��2�v�h�]�׾�6�^��}оV \���>oW&���нEl?wF��	�m�M�?�G��I?	Z\�t�
����hX�?\q�?* �?���?�C?݋�>�Qk����?���>��!�G���[w�=�=�>,ۿWm���ؿ������F���Q~��?2�>�}�U�
��hx?�޾~!�?�`>?�I�>��7����>/HI?V���G�L��ei��O)?�7�?/��>�@?��>��X��C���Ծ�L�?���\����՛��N?���?e� <X�>�"��Tҿ_ǽ�<�>�����td��?0���>�I��@�>L?O|>��j��>Ae۾���=����z迕ۧ����X
@K���!c������tZ>T��&/<���罉#@U��>�U;�^����>�뾩��>�a?�8{�xx������2�9�ؾ�T?�>����aY~?�N]?�����>>��=����훾)Q>��j?��5�,ɴ�����md�?@�>ђ�?�$ݾ�kT=�Z�>�%S�S4?+_�?��6?��M���[?mwM?ES��r�> J�?"��??Lc
?���8T�>������L�8^���ܷ����>�D?���>>ߍ��w�?����n?�M��mو�x�{���D?u����a�E�?�?��ſ��? K��1Š>�?�?�|Ǿ#�?���?.S��j�9���3��������?m.��w�>H"������$@fM�>�v[�)��;�@F,"?�묽ȟ��)n@+x�?J�>�F.�T���P�P�[?�s(���p��lT�lly�T�0��X�?�s�=v��Lʇ�&4�?)�>ܗ�ߏ޾E?"��>c&��o��?���c�t?���>
`���=�6፿��>̱��G�徰���վR�>����>��̾�bv?O�?_������� ��XI@>R�?��B�^C���ї?��I>�O�����_}���e??q�^g���!?�7?��a�"E=_�Q��?b�?r=?�nu]�^��=DB8�@<�o�?D*? �?�tI?�x@��?�b��r�I���O>��?�;zGw?� �Ӷ�>��B�u���Q�)���R#?U_?�eL?�;�Ԝ�+e�w�!�C�?ZZ�>��>���rV?G���bj����>h�`> @8�.�6��о[�A�΁�q����? �ɾ�Y���C>G <�\�<Q�f��>�><��:�H��H��?��%?�
��}���*�?��,��Gܾ�鉿۽�=Fk'?.R�>�>w?��>��M?�臿�.����>VO>;]Ǿ<̓���>5��>�5d�k������c�~��n1>X')>2X�>O����c�KV	�H�#��=�>�z�?���=�X��g=��	�ʽ�e�=�W7?��:� 6�z�
��}{���Ҿ��U�h����~��,2<%���=�p��/7O�Ƿ��-�=�V�>sǘ��0��5�N���F@�4?�N
=��>� �?*��>p�^?��><�-?���?��?��پ����C}��7�O���g��>v;?ˢ�<�I>�ۯ?&�%?EM���z<��<��?/��ܺ�?}B�>��>��ؽ�}B�1�-��>��=d���p�ؿp,�>��1�eN=槏��g&����=_��>�>�@���^��? ٺ������_��>�8��,� Nv�]"��|�> ����E��2�<	��?d�?�҉=&d&���I>E��>OOS?8�>d->M-ǽ��?� �>�@(>�����>2dվ���:��>�L��"�O@J?Ӆ�>�载
�?��?���N!<M�>ǆ
?@�?��.��g��xw�#���q@��Ⱦ�?�#���m����?�?x?��U>�����=��"9���	?��>�|0�(0�=Wn?�r�?�D���Ѿ��P�O�>.`�>�M?o/�-f��|(=D�>���������ۜ�?�M?�?�k?+^h�mϒ���=>]��\�Q�K
�=s�K���o��:?��ʿI�=c���*M���C����-�~"�7[�?��y?2�D?��[Ws?�S�Z�V?�F(�j&�����_�?3����_�J��?�t�?>��%��?��?�\������D�?4�.?���?���:��?(�?�P�?}f��z�c�Vb3?�1�?��&?��7?1C����>$�>��`>q9��a�
�?��?}��>�h¿�2�����Hx�I�n>��W���e?eya��?P2(�pO?q�T�5�@W��?Z��)���?�ry:�ѽ�f%�^v�?Q_����>�����y�?}ړ?2F>r�?6��?��!���?>�	>���?���?�UO?0�G>��6�?�@�?
���Љ%��|?wb�{�>��T���P>X�>���?����ľ�X��C�=?�����~�> n�E>羓��>�k?��>]��DP��mPj?d�>�y>��%g>п��*�F(R?���=(����=��3?�l�>P�?��ƻs�?M��>M뾊�>�7>r��<N�+?.ý�nP��A�K�:��{>�(>>�8&�b��w�A-�?+�n�̯���]澹��?���?���?+��?.g3@&.�>���=�&�=�徭ǿ-?�>�~u����<o��=�|)� !����><d*>����Հ��*�P@r��>+�I?�Ⱦ���?"y*?w)f�Yve�D�?��j?s*8�X�O�}�p>%~�?�� ?�ӽg~���[h@��;��ſ�6G��@w[?a�;��o��H5@D7d?F�7>��s���?i@�=�?�	�?�"?K�g> ��>Ht)��z�%�/�T?�i��Rh�i�>�W���E?�m羝����(��C ���?��?�(��y����,��4G?ɬ�?�b=qt�;]��?�o?J9���Ռ?� �?��>���>r�>�t�<1' ��-�?8GE�z��@��[�����>�1�?�Ǿ}��Jl�(����0j>ր�>v�4��P����?���>��?��Y��d���I��0���������9H?�0�i�;��؁��vJ?�|C?=j�?<�ǿY�(>��n?�.�>6�ȾśN�
�z3/��h�?�z>��0�ނ�	l�?SG��}"?���T-���>("���0�]@?�C�>;��=H@��׹ͽ��۽�a��]���o㡾Ƅ>��>X�ľ妖?E��?Bۭ��?�:>��q?��>�~?�2�?���?��[?1n3?EO�+����>��)?4�.UR?p��?\z�=8N���>��<>�4?[G�?-ع?���>�N?���>bS�?��9>\�6?u�L����n�A��=	>�\o��H�z�C�DGy�����a��P�>�P��:�Ŀ�g?үe��{�??�>2f�>���RW�?�������>ܜ6��Â?ͨ���9����M ľ�b�a-����ܾ^R�?fR�?Ԓ�>m���*�=Զν��1>��>?�Lp?��Q?O;���خ=����A�Z?]��>�l��gQ�z0?�z8��d-�㠿w��>����ؾ�h��.��Yw`??V�?J�S?s �?��m�MR�a��:�>�G=�$4>@�[>�u?͆�>H�i?�}}=��#����?+ Y?�8c������Å@-���=q����3�?�t,��#��2:����@���b���:n1�/�]k)?'.���G=7�b?yZ�^>�E^>򘑾���V?P�>(�F��1L>��=J�����>��?ըK?մ�u��w
>XǷ>�Bվ~��>�ȯ���ھ(y��]��8m�<�S���_���Ҿ��Ͷ��p� ?�.�>C)?�(g<J��>���><�|���?<�>d�>I�?A�'?nW�>�..?DN�H|���G[�jIV?��<���>]�!��3y9J��w|]>����@2�HԾj�,��&��y���-�R�O隿/۾���>O�����?6��%8�>G����gp>�;����)?��!?&�?f�H>�b�3q����=�e?we.�������� �>I���s�^	� ?��?�O�B�#�J�>}�ǿ�����¼�7���s]���J>T(?�2���3�>ĵ��9�L>K��?1?�?��?�R�L�򽸪�� ?O~߾�9��=���;�����D���ѿ�l�~)������{,�>?>�}2?���> {�=�>!Ug�Y1k��Q�>�+Ӽ�Kt������B=��z� q���:T�(ou�6#���~�Ѓ*?��!���Ǿ�U�8Ͼ�j�>��J>�����龠7&���)?��ľ�q~>�b�>�>c�=	?�����V���}�>�T�&��K���/�/?��>�w�>�}r?�1�>��h>�Ǿ7*�@<�~E�~��>��=Q�,>�o�Gn?���>Nl?>�9�F�=�����v�?\V?�Ͼ,�=Y{��T�w�$/%?��?ܑ�>W9���p?�𻽍K��~T��?��v\�u X��ۛ���='��=�+t�^�1>�6>(�=q������>��'?�u?������>����� ~=�}?y��>L�?���>/�>&s>��>�aX�.fB>-?�����ׄ>ा1
�<��<?��O���f�)%(>y[��11?=~#�LP��9i��?m��_꫾l�>��3?tp�>ݞN�m�>if"?���>;�#?k,?�5?Ƌv>�.�>�Y������Ax�Q��
� �.E�?k�/���=��>N�??�0b��5�>	5�=o��e�9J��J�7��>M�����>P
�q� ��U��O�O����>�?��zF�.ڻ�ٕ�+j�G6��.�<L�?۟(����=oB����^>������ �>� �>���?�YU?J�>�%(>��i?�Z ��S�>0X���>~0B?):۾�得�������F �PǾP���U=?vrz?��>��N��_z>��?�>��}�z�?���=q�B>��	��S�^�>�V?V����0>�ľ�5�>���>�v��_>�G>��>l}�-�>;�?r�?#��>+� ?[7?�?H;��>z�J>��=m���`]�o:Ⱦ�P�Y��x���Y+���8�U��>'��=�E���循�Q��$����>��z�ȶa��"���ů�p.?�������j"�jlG?X�#=j�z>���>鲨��P���V?��=>��ν��)>�����=w���<	�B�F�Hס>�?�H?��>N<T?�ܗ�t�������$����c>y�>�>ԾJ4�8�$��I�>Z�����>k�>u�=:��=�Z>:��=,�<��O�A7Ⱦ&�꾸�0=�%,�p����?6E?!=a��%���v���2�=*9/?L�?԰?�k�=��%���<�e>��>�#L>qx�M͇>ġ�>=\6���7��Z(�w���󨾛[�W�����A�z��@�=�/��Ȁ>>{>5̽�0?i\>3��:��y�\�H�V����^0��O���f7>�e?��>?�.�NxQ=Җ�>�Q?aRj?��A?T�j?�;5=p�;~�ɾ�a�I}�;�|?�2�>���> �o�����9F?�s��0�=��?�AO?N|J�T��5�4��2y���㾂O>lF!��齻�����?�x���lO�I�p�6��>��1� ���IU� ��>D�k>>�þ� ��>�~0=�ͽ��>� �>�
u>+l_�gp�n�>a೽�G�B��>��K?ʖc?�զ�Ȯ�>���>�x2�ڙL��V�=\79��^�j�>Z:>C.�����?Nn��&�*>�Η>�s?ߢ�>��2?�2�?[%%>��?�I�%-H=�%2?��&?*�?��>�Ӿ?�������6�>�k����L���=�-��Ȼ?jՄ���X[�?���=n��=�P\>>Ȗ����>-��>�x�?�M,?U�?_q�=���><���z?���=�_��ϾAGv=I����~�bA=�O�=R7�>��e?�J8?Y|?��5?g������߇��G?���R��މ<?!��=$���4�Ye�>�gS���?���>!⻽⥛���׾Y�>.%C>]5	>�)I?�����3��N�;�$%?����i����T�Ļ??'�W>9�����?�JZ?����>�*	�n��>YU��*�����Dy���Ⱦ&>���>�e??̍=�R��Z�||����>��?h��F̋�d�t>�|
?�R�=�1i?Tn�?�Gh>�I�>�m�>"!�<ݾ�ET�\���>�뽋� ?,L��~<�>�>��RBm?ʃ����?\�>>�׽����O��W>BF|>��>q&J?�|$?�>�l?}��?��]?�{�>^(=�w?9)Z?��P=-Ѝ={Vg?sK?�w��q�]���\a'?Hǎ��럾-�>�"?S!9���>MĖ>�ݢ?�O5�%�=��j���>s)\��uy=0>P��э���)f=
4?j�>���'�Q>�ޅ?��j>�2Ⱦ,h����?�b����>��־!
�ܸ�>�3?i��=̡�|��=���>�?t?��꾎b�����?�ぽ���<z~0�oC�=B%�->?f˾��>/��>m\�>v�f��=���T���<->��>j?[Q�?-�?ll�Y)�3�>&=��K?�޼<�N�>�{O�0��>E��>c�������sƹ��������.X�3�����N&�;�+$<F
뾍Q%� i,>�I)>�=>��>;�=��j�G&��I<��%����}��U<��>��8?%���uz�}xm�bU�?3�~�4|¾X �	,?�T���>o)� Cq?�����>ʫ�hD�=�n�>R#���2�r��=�xý�˝=x��Xڶ>��������۾@�
?dR�=���?n8Q�񬨾&�=���>�2{�`���&���>���=�=L?W�n�k���亡�ݾ��=B��>�� ?&9���5����>�L��I�����o�5�?�I�>.�?�[���'�Լ�l�=���=A�>�f	��u��@�n<��?�{�ȿ��R�v?ڐ>�Q�>#K����`?�8?������?.d� [��5$�]hF���>��>�`��C�>����$?�d�=��?�y??�)?��Y?���> ?	��F�?,�<���=G�z>{
_?q+��ߺ޾F�?R�>a�2�R�
�B!?fFA����J<��� ��!��!ܾƥ/��A+>U��"�嶪�7;>��?�
>3˾�>��{����=�ͪ��87�1K ��aܽ�T3�5�O�!?����P�#�ɂR?�Z ���E�=��>��?�'�>�t�?��w?��?���>�2?.��='���ps��Q0?� H��v��O9$?�>�1뾢�k�և��Y�>ç�>�y�>ϥݽ���en>*�	��qؾރ���(�>��`�y�>Х��L��>M�̾|඾�g]�HJT>��<ׯн�>54w?�?��>
����Y>>�?�z�=�y� 8��?��=>�<��ƾ�vӽ�B$�>J~>]C=���>��O[9?9]G>J��>�8>��?��?>�@>�����>u~?X�&?6�C?�t�>�H?��J>QL>� ��bH>������J�$?/�>���=��>6z��^r�>�6��Oz�o��T|?_/�>�0��[q�\Ŕ>��!=��=������<?�ǂ��&�>(xM��{�=\� >�� �s��=ȇ�~i�5#���8*�`��3�W�QqD�Ask�]X�=��<t��;+k�:S��=�>N��=�X|<��
>�l�=�ɍ=�{e��=`=�fx=���=zE�v;w���p��.���[��7=��m\���K,>���;�P�� ����Z>iK<��0��D����=s�>�kb>��
>�p�>PH��]���1��� `=X�=�7<��j����=�P>>���W�Q�=h="v��U���w��0�v�j �8�@�f�E�˗�=��=�?V�~�<�n=YNf=Jf:���f=��=
p>�i[>T�M>m��=2->`j�<`G��l�;�/z=�J����[��n=Q�.>�KM<��=����:�k=�d=�ꬰ='"�=��y�?:=G��=W4k=U��� Iټƭ�=�ݝ>ﾮ>�B�>��>�Kֽ6��Rͽ:��<�Z���8���'�=I�L�_����� ����1��*~��t���>�"�>K�l>&�=>A��=�U;-��<�=�mg�\��m��5B'=�[�=���<� -��g(=���=9|�=�3=���=����w�]�Hr�=�:ּ�ټR��=�O�=;��=���<D(M=��)��G$����d�(�p�h=��x=\�0�XEA��?�=}�>>c�>�y���틼���=�p> �׽�+��ν����)�����(ӝ����=�X�F
��P"���P$/��Zo=K�[=U�=MJ�g0=�|K���<�a�[�=�v�=n"=�Tս�F=r�=e��=m��<��_���L�$vL��kp�P����Ӫ�-�l��7d����=3��;�����ݡ=@�={��=��߽�ꝼJ=���<�NսRZB>��I=-V>R�=��<>��ż?>��	Ȕ�"e>{��+������;>$�/�!Κ=A>���*�<�}:K�g<�>=96�,f��MP�y#�>���3���KEQ�)��=92�<et�*Ȇ=.�v>�ҝ=�Y�=��Y=3<}>I�9<w�2�+�g��<�=��?���C�+�l�f>��b�����6<�0?>�L4��w�=^��=��)>��0�v�s=�1=�v�=�G2��W1<Yv�<��=$�i��G�$*���ݽCF��D�W�K���{Қ�)���N����
;�l�s����y�<��=}�C���=�:�<��ļ��V�0�t=�^�=u}�#(>��>|C�<1����!�<�i�`27���`M������9�����^���	�eg�=�>�=4��=ZM� �=m	>L��9V-�X�3mv=��=�l��A�y��t;��n�&J
>˭=@�<�j3>��<l�ٽ��-��<>6��! ��
I��>��=-�&�w E�h�=�N=��:=��;=�t>Ҏ����r��͏=vW��h=�H�<�7�=�<�|�����J�k��q�e=� =�+t=�%>3�X��:^���Z�>/$��I��W��v�=��=+J �\4^=��>۔%����ԛͽ���*�=����>=6(�=`�
=�'Z��½C�=a�B>�Л>Jld>�>ԫ]:�&�y��*�C�:��<f�ǽx�ܼ��=����͏����@=��>�W�>R�d>��G>@>0�v=�B�=��?>�:�=��{h���">hu�=	��=����<�Aq>Ӫ:>iV>�+$>���=nk�=o�=ΰ<��=K�˼�Z������D�=l��<��=�׃�a���x%���t��H�h�x�|W�̟���a� ����|��^�Խ܌t�U�_��Z��S���᠁�?�=���<0+���I��3���C��B=6�5�������=�PμLy��Dl���໋!=��s��3��.^o���C�������:=�/=�F�=K�<Z�/���=�s໮>�k����
�<�> >�����(��]��\Uy�Gp��9P>%��=��<��=D|>Mo��lR���	=2�>K��Ш���D<( M>�­;B�=�m�=eb>�փ=�6�����=�#�=��`�н��J����=
Ů��V��>�/<Il>�D>q^%>�G�=�D��tz �"���P�=����.;�(�Yf�=�&F��%T�N����L�=a�i>N�>h��>��\>�n��	 ���u�;
�����30=�$�7��9�k�d�,��,I=5:��Q5���T��2Q��e���']ؽ��ڽ3�<𽳑��2�o=m��=�.��^�<.&=S�=?�"�V!�5ʍ�ﻘ�<�c����Ǽ�Gw�r�J��m����=P��ѳ�=���(}ݻ�bսU2�=`�^>�h�>T<>�l >q���)��,��i������{�&ا��'���5��<�s��������=���������>�>>.� ���>e�<��D��D�A�>�%��{I��ԓ�WC'=9a�=��;��x���@>̃	��J�;l��k �=&��G}<��3=k3��̲:�ܜP�@�=s,�=�?��s#�-
����U=��<==J��<,?�=�5�<{Q𼃒�;��U�+�<�Ӽ������e����8����bS	<��=�>�<�L!�-�r=U�9=�%�=A�R�ߺ$
�=r=~?�{,�R��սԦ8�bA>�g>�ݼ=�9�>J�7>V�X>c�d>��@>Ȫ5>?
z>y6�>��c<*�>A�;>UJ>�>��ʽ��>��>'M>_�����>.�="��=X�@��=x��=�>a����󴽦s��_���)�b��.�ǽl�½�g�<��<=Tw�=55��ni�=��=`~�=�/C�HL�隂����E���w�J������u<��;��D=0�+=	��<�F��4cG=���=�>~9M=i������J��n��U�ül��;��6��O=�4Լ�I]��s�<d4�Ts�<G�6<F����/=�l�>_Q>,�>4-h>�޻:4�?=��:�)���n=>��=.�j�>��>�19>���=��4�=r�ջ}M;�4o���,��;��솾
�<��=I��r/�����=$�'>%�=ϙ��,=��>���=V��%y�{�/<kg4�Qu=�5g����=4�=��=�ʃ�j̿=:�>P\>"���q�hR�)q>© >	��=�V=M{�=
�g�TU'�3�m;&rμ�n�����I���D)�=K	=��;�X<�<L�i�e=�<vb|=�>��{�=�²=*W(=B�#�ƌ���df=�_>�Ӌ�a�7�G���v�,!���{�=�N��U�=n���~�m=�V)>�g�Jٽ�����t>j?�=>H��v�ʽ������q=��<х�����=��=�VR=Pn�=\�=2�>���=XT�<��>�E�>sD�>v�>%�>lk��}�#��'�l��=��*�U���s�;�#>���/�=����s�y=釗>ݓ�>���>F2e>
`���=�U<>��"��=�I">��>ޙ"�{A=��<~1����*�_����c��L��84���n�m���w�����=�Ö=��<��Y�oo�=!�=���=�u�;\:ѽ��>�:��=<�o<�z�9�RN���5<���+*=�����9Q��lM=��J�~h\�L
��_=�s�>|�><Z�>㙓>$�*>sͳ=r�>��=1>~&�i%��ƪ<W#Z>6�����J�
��>���D�˼���v譽��=�{��Oh����=D��;z�;�f����=G<�}Z=�ތ�zd�҃�T!��������b�֢����*��G�za?=.�y<\:�2A�=�p>��=�)���9���h�yT^����m��/�G�����G���Q��=��!�"�(�F�z��2�=/<@�=b�U�{n���<��<�~ >��=D�A>�1>D�>�6�=*��H��_�>e �=Uf=��\;K>���T�z=�)��^�IIսF���P��i�2*�b��	���!U=��Ƚ�V ��T>�9[{>� �=���=�g�X|��V&���hB?.���?ξ^���>�ɾz�����H����q>
 �?jV��I�>��p�qw�?F�?t�?�y?��I>��?es|������J�{�iX羘\ >[.�>����r�M��p�'?:�1����Y
����d={D�81/?�:?O�X����$D��?�/�>���y"?߈ ?T� ���<>�wo>R�>`�@>	��������]�?H�>�$?W��(>S��~���@�߹7��"�ց��D#���=�Фʾ�L��ii�>W����>/�о�2M?��Z=�(�>��]? �_��>xp<�w>1�7?I�<�{A���j���>�'ڽ�dz��?��绠>u�?`þ�V>e��>�oO��?h0M�����-&?��������h�>� �>��d��پ�FT��BD?J&?�q?�?�R���"D��r���t���>�.������A羨�*��ߍ��.���Xܾk�ѿ<��ë:�8s#����<�8�w��>�J�U�ݾ�Tྗ9��\=Qdy��)i���oc����=���=�χK�
DP�Dˮ�3������?zn���ER=S�G>:Un���D=~	>���>a)�>��?�y}��\�?_|�$�@?-�l=�L)���>�&�>X?�=/��1M���>�>?ي"�Lƛ��=�>���=ߴB�/�1>��վ2�����J=?��=�+?
�??��>�v��Ο?%)�=tK�>�U
?Z6��{ќ��5>� E�F���@?
u�>`�>+.˽���>����#Y�!>�?E'�>ܥ�?2{�"� �A�S�&N�~�;���l����#����>�F
��x?n�X�to>V���Tf?h7s����>�c�>.B��˽?�o�P�>g�>���>��>d��<03�>6r7��d�~'�r���_��>tʝ>f� ��E>~�=΂�>P4�O�k��>c��>�?�'��v�i?�����>)�7>�F;?�T��.y)�%B��:��?5@>3�=?
�=*�?t�����r���?0s\:�%?�Y=��TR��N�>�߂��B�=�/>���}�^��l�?���?ֈ?´�:Ѿ=V)?n/>�tM��ȉ���?�k�>�U��踿��?h�ֽhW��BM�,Q�>I�4�=�?>2)�,�>�7 ?�[��B?��S��>�P�⢅>ro�>p�P�^��<;��h�Z?]&;?��ʽAާ�~ꜿ�0�(��� I�ǽ˽rK�c�����i�+��p��8�D��?��(�蜡=5y���:ͽ�?��	>׆ᾄ֞�{׽�.#���`����?�@? I���>{(6����=���=��ri����:=7@�=0s1��`���ޏ>B\�(��x/��o?=�*?e�b?ொ?I�d?�����5��C>	˵�{�����P��㾎l�>>�l���2�~�߾P&>fļ=���'�=X>�6�1�դ��4QE>2{=R�b�EP��� �|���!6��`�>���,��>ȦA�l��=2^�>�L�@�A?�é>�-�>�-\> 
?��˾yLL?�w$>��޼�]����Z��N=�Q���ž�\��,�X��d��}�6����݄>���>��ݽ
��>����_�<9�U>�*=�=)S���M��聿��Y��f������1_�<5��>"S����E�I����G�<9}?��?�Y�=�FN>4�ܼ8�=^���NG4>��,?%��������?���H�2�c����.��`?/�ᾢ�ԾJ>5��n�Pq=�l�����A��ɰ>^?_��>1 �zA>�{?�![>�<���^���k>�ś?��s=%>?9�?� �n5?�C�=����Og�1|w?4�?Z?H�=�09˾��C�32�B�?��>��ȶ>�; �(�� $��x�=z��=2�?���������=f߽>E�?(��>�e�=�U���u�����[��=32}��%��\>�R��%���N����h?}6A��s��a�>�Y� ��(�M�KT�>�t|��a���ȥ�կQ?�j�>��n��7��*p?���>[�R�[0?���>�\����?�g˕�x�x>TR�=�E>7p�=����3�׾� ���V�m����H>�!1��z.?�����fk>���>����??�:�>�9=%���s?��(?�l�?p�B��QG�֪z��!K��Gi?h�?��5?x)J����?B�>�X?ۼ�?3)�>�4?K7g<(�S�
�����?��e>Kc�?����w�=X<?��>�E��7-=�z?�3v?Z�?��>e]> �=�j�>�V8?�0�?�i"?�3_�ݞ���V׽%���b�����=�A��~�$���<���*����u⊿�td?�O�����w����[ཿs��2?�;F��">QPE��rx�:��>�����?<�?�>g��>�c���1�<#�;>
��?ߤ���^?Tv�=�r?߱�z�>-6��]���Z4�K���� ?<;�����~Q(���T<0�+��[?��9>��[;��?δi� �1?�qX>�������;�>�Е?㿡?d����Ǿ(*�Ҋ/��h�<,��?U�?�
>?��5>������D�P?<��>P��?��J=�ر;������o�z�S(?�]+?��N?.��>}?M�?��>�?1�v?��T?NO�?a?�
??�?o�P?SWM? ����?����	�?0�i���=c�)?A\�=�}<�p� 2n?�kQ?R��������<&��P����=Vr���.��q׾9�>aۮ=�&�H/<>}ۚ>��x>�i�������	=7Tg������:?��>)"�>r��~i+?��>� �2A2?����=�C;?Շ��PR�p;?h3<�tM�>:���k�DZ��z�Y�D>3���`�=���>`\W?�_
�
貿㵐� �>���?q��>��?�-����?�S>�]�>Q?>�7�>%3��sĢ�� �?!4(?=0I?n%¾p��d#����ξ�7�+Z�>؝>��Ͼ͕ҽ]�Z�{�y?��>�?���>/-h>�i/��>>�s#?�W�>��>�2Ѿs;��4�A>�i�>��.?"jǾ0�!?媋���>���%����?v�s<O�E����K?�E?Pu��7���p��3��?�٘�<o���T� �=�C�_|���4��U����?��N�ۡQ?w�Z�u$=�ʽ?)?�v?�Ol��a
?�^o> �9��-w�\4���� ?��>*���=�S�=�� >��"���?3�þ�g�>N�R����b`7��b���(���f�rF�>����uo�x�(�#��>-���\�> 
����ϕ߾b�վ
諭?{������^'+���>+v�=��b�HžŴ�>XM&?��>[h>���?f�2��% ;��?����(��!��=c�?L�2=��x?e)۾��R>��_�c�>��|?�T�TB?"(�?��]��0w?%=�=�k5��c��Ȼ�?���?�E-?�p)�"��������2o�lP>|4?p�M?V �>I�>sz�?�eL?wi�n�Q?��<^Z�>��?����qj; `?�V�=Qnz���>4Ӿ�'������N܁�:���hx>+V?m�"�^ ���տ*
?Qk?|@?���=���>ാ���X�?[84?	/'?�W>/�>b��o/K��r����v>p�#>������f�EB�>b�8���߭?�����&�>aّ�O����h=����9���m>^3��#i�>��0��|���������F?�"�l4>�ټ��%�m
�!%��	�G??�J<���?��]?���H�>>>y�?�z�>�'_�΃�=�?�H^>KYb>�?�VU?��ɾ��� !�>���>����1Ͼ��%�:��>�O>?�?�\�?�?�\�?�GP>�e��<c<�8�X�+?v��'=?�>?~%?��?�'?��?Uy��S+���������a>�$����%���>8?|?Puǿ\G�P�?WĈ?�/��	�k��=m���Ί�<(�S>��=s��a����<"RW�Ow���U���:��>�LL=@�k=��/<0�">i�&>�b>TRٻ��=<��=��B�v=\s�=3$B=r1��Xo��82{�f�8�u!9�Vn���Q�S�����=���\�Ƚ��=��>�j�����Ч@�Q�+>d>"q@>#0>�x�>p�?��3�g����H�qm>�=�t�=?�A���=t�=Vs�=	�R�w���pT=�?B=�`;�nʽ��H�ۤ�71]���u�\�'&�<q�=���O�｜	�=R��=OϽ�� =��=��=:7d>=�=��<��*>�=q5���$�$�-�[d������a����<��g>�W��@��g�=t�6<[�ȽJ|�>F�=��.��z�7]u����=]䀽�����^{�Ѱ���>��)>��>61>�Q��v��E}��M]=����e��匾ȧ�=O�l�y��;��n��Ep���?��t�O�^�$0�>�L>LI�=-�>�k�< ��<�{�;d~���Z⽅����
�<�.@=����HX�KG=Pg�=�X�=��=xϑ>І�=��=e�>��=U=S���b>��P=��>e�/>m*[>��>�g=�Q*��yq��Y��)|���0V=lR=� =}��v�=��=�d+>�m��h"���<Ǡ,��ܐ�sjb�j�O��6��汾,>H� �]���h��F=�}��m��=5��<l��8�<�R=4�O������=�N�=u��=v�ǽZ?>�N�=a_�=��|O�=��=�)�=�c�ȣu��v_�
�t�������`D4�QZB�l�}�d{Ž��6=��*�%�����<*��=M��;P��r$罢�==���d�.�">�(>F�=u�~>��h>ʋ	<�q�=��Z;��j=T�񽚶N�Bp��s�>5����I�����A>��L>�E>�]�>�n�=�ls=o=j��>f=����1�����>��
>��G<���=��>�#>Y��=Ʊ$=�)e>�D9�������=洖>_"鼟���
��ݷ�>��w���ܼ�6��� >,@����>�7s>��?>#��a�=�혽3_>{ѐ����=�\�=�9=��͹x�㖾�n׼2�����y�ٷ�3���/s��q��=$�m�}�<�I�0L�!������=�����B=k�R�>��<�>m�q<��7�q�g�j�����_Tɽ�G� �*��]B�KƝ��JӾi������,��1��=��=��3>캔>�c���*>��F>4h�>�nV���)>)^�=U->~i3��������7=�>��x=#��=��H>S��</q�H�,=/]>��:m�W���Q���=�\(>���9�G=��,>���=�LY>䐔>2�k>��5<]a�=�� =���=���ƕ=�;���=��r���:���G���ֵ�=Ժ�;�%��I�=��=���߽IƽO�g=��������x��y���#>�)>���=���>Sm<�:��q��9����콴�<bt��'�=�{�<H�f=9�=X,�����>y"a>(R>>�`>�î��w��l ��t};��T��e<�!�� � >
��<�P�=z�l=�(�=�:�>���>W�>Yt�>cۧ=�ˤ����C�=�� =���-�K��>���<J(��`D�hM<��>,iq>ր>{t>��)>��>)�7>�~M<�R=4wq=uNؼ�D�<��=���<���;F�N�j� �e�#�ܦ{�({���O��/1�.�N��f�s3�!k0� Pn���ȽmvK>,��=��n=��B�S��=�N��P��<�Eؾ���_2(=j>�]��s<	��=6X	=_�<Ŀ4�PI��x��!f#�����rY�:����^��+=��F>��S>'㎼ë=rl�<}AE<8��|0�Kv<����$�=�U�޺뽿ƽ��X���,>��<�㼼<�<�P&>����LG���0�&>E����m�wlg����>H>2�=��h>%�>�Ć:z�y~*=ݒ�=ˍ��o<��4P>{缽:��j����>�9:>/��=")>VH�2���I7��O>|����ۻ�Y�=�;i>AWR�%)j�,QĻ��=�{o>g�i>K`>4#[>�q=z:{>�EO>���=�]�=z}R>�D�=��Ļ{S�<�ԃ��*=�;��4�-��2��E�]O"=�p=1$=�X,�Lr�<1��=_�=��u<٧!>>��="��:+�^�;=qi�CĽ<�F=X@F�Ľ��ɼB�[=Y�:����=R��;v��=�I�=B��=t>�%�>�)�>j��>S?>UZA��gp�֬�����1����^��#+;�괽Á�=��>nP3=�BA�z4�=0��=5z�j7�����>g�d>JG/>��>�1�=<Wa= Z�<Yh)>����Z�<-���$>/�=��E����=5<[>�uU�ݽ$=�h
>��)={м��CF=1Ġ�W�*>z?�=�Ɋ;
?�=�֟�u"J����ҽ��>#TL>;W>��l=�:>�R>��G<��U=J�	=�
>'�>n}=w=��｟��Q��@v�>P�'>2��=W�?�q">Ԏ>Χ�=�Z]� &>���=��=|�]�:��<�PC=��Ң��>
�3>�pg>r#�=銚>�_�>&�>~rk>Rb�>��>_� >���=қ>)Rg>�]>�ҫ=� ����=Ǩ'=^�B>�!T�_.
>9�=5g(>��Q��]E>���Dd�=^]�a�����=T���d������{��[D����3Ɛ��ֽ�a����s=��3>F�;��G�������	�P�]珻�|��ә�:�8���8!���<��=rzn<O6����\�v�F�^=*�:�Ҭ������>���l�<�h��uE����<{,���&��zp=��ďbu��_f�;�o<�|w>�r>�ds>�>Xy�<f���� ���L��v<E��=�B=�I�&�n�����=���	�����E�`�Ň��+7�I����n)���(G����<�%�=BB���D�=���=1F;�c [���<����ٽ����+=�1�=H�>�A�t��=��[= ��>����e��=:I>�=>����]h��	lF��(<=��=ge=?<�=��4>��㼨W�:�Ͻ���
��<D���J����=g��=a��=�D��y-:���*=��>=�g>���+��="�=���=�՘�;��<�Tb���G=^���<�U�X�>Sq�f�J��1e�%��=�
>����-� =�*�v��=�G�3
>�A��|S9�y����
�̛/�R�e��ER=��*���ǽ���=�=�<R=��<{��=��e<� R=�3�=Gw'=߷>��>��>���>�7e�������罗���T������Z7��~h=<�������`<�UB=DЧ>QL�>I��>W�n>�>'��:�+;��-�B�V=�[>M8>�&k�`I�<��8<)Ț���=�]���~'����0,���}S=)�#<�d4� ��=��j>���=�6&>�8��|�=J%>��/>�=A<K�̼zȚ����<��P����&��:����ؽ�_/</
�=Eh�;�Y���S���6=�\> y>�&a>�u>��<��|=:��>�,�=�#��� �����T^��� ����Q�=�eT�T�k���L�� �=o�=�W�=�B���ڽ`DF��}��[�j�&��q���J�������;
�������)����S9��7�iR����s�� =�%>$M<d���s�=�[8>Zxu>���=D�����<ٽd<C=oA^���T�q��z�������̭<�Iv<��9��u����"=�>��="��PA�!��GL]���X>Ɋ9>~��=�A�>L�x>J`=��=��2=L��=��g�����'��u��=�t�9L���%�$�?=}W��6�^����=5m���p��q�T�Y�Z>o��Ȋa��S�C�>
�T=?��<ͺ���=�m>[r>��=ka=����<�c�=.pQ<x�;~xؼ���=�s�=iV�����=�>�Bg��>$�==\@=ݑ=93P=�=8�W���;^�=:N+�l��lsf��$l�nU�kqI�[��=�ސ�K������=0�4=��������t>���*��<��l=r#>��>��>�ge>Fx>�L�����T�=�����=f��=��?<�c��1/>�o=��>�췽��=o�w��#|=3��a���`��1ǽwl ��))��W��tj���=72'�"@���|=�A�=qT<�9s1=��;O�=xG>T��=��	>�->AR�<@<���Y�M�<=s�O���e������<�Rp=���1j;o��=���k��I5)�#0�Aڵ�h˽���U�7x���4�{�H��oy�����A>��!>�(P>B]><�*�r[����!��(���ü-�����V��b�@��I�AJO��U���ս����
}��0(�&e>a��=2\'>.�>�϶=G��<��:<�Iּ_s�=8xC;f2���^�]uh=� A��.d�R��*�=&�2>z@J>�>v��=��t=5��<F}=ľ�;��:=G6�<���=�r:>�Һ=
��=��>��:��&���ѽ��V�)�z= ��=16��M���.�=���<>�>��Z�#g�=�=�>��S|8���0�])N�x�ҽ'b�Q-=����c�=ܲ���V;��:�=O�>��,�RM�=' =��>��;��?<������6=�?����=;������yb"�Y��=�<b%e����A�k���w�������zͽ�<�g��r*��mc��v<p�=ŝ�Cq��nW-=w�=(c��S`=B���S�<�)�mdp>�0><F]>�*U>fy>�@=��=��b��Ze>%�$��?+�v����^>V�C={�=���<m]>v�=�ϧ���y>���=����K��>�>zVK���<m'<�N�i>h"#�Y$�=�0=ƃ>�a8>�]L>Y{�=u��>�]�<�+=����lQ>(��9p��Ce�<#�,>'�C��ӛ=!�=�+W>H�s��=I�a>��X>q�ѽ��2=�]=� �=(T��W���;>MEb<m,�����˽8��aU2T���@�'Ӆ���G���]� X��5�A=��<�^ ?<H�=ԫ,>I�<S=yNl<������=��=�B=Rͽ�
<�n�Z�K�@�^�<��/�a�ӽ�<��H�t�V]��ji�[�s��	0�� > ��=�t>%��H��=�g�=�E�=ڜ�.��<˖�=��X=xh{�v-@<����������=�t�<��*<+~>��2=�N	�D��6A�=�A-�yN�<t���0 >�t=�I�=O�8=^(>��
>;`>?X>1�>�L(��B�;S�=l��=���>���j��O�=�M9�&����0� ���$�=��=i�<�}�=��z������(n�=ba���r�������'+%>?:�=�@�=/~>C�}=��M=^PX�����n9��������G���<�=�rƽy��<�C�;��E>��*>F��>���>��
�v=b=�Qｹ�<��T�^฽\����� =�e,=�n�>��<J�{=g�r>7XF>�ly>6�>)��=n�P=�*���1=�e=�c����҇�}��</���7���0��	L>�>ڬ�=q��=1A�,f=;e>��V<�&=�)�=E��<�i����=S]�=�B���*�����\m1�_5d��,���k�Z6��[�ƾ����
��C�4�^�i�������ۜ���>��w(Ӿ�}���-�V�x��n���<oy.=�>eyM<u`���$=H=h����ͽ��'>��4<��5=��_�������T��D�)t���6���>q6�;�#	=��=R��=h�=bн<ln1>��i=�E�=��V�cd��D�9po��PT>���n=�l�=V~�=�	/�-���P�;pJ�=�}���p�&<b=�;:>�j�=U��=��P>�>��;o�M:�6�	}S<��۽�����e�^l=���Z7�y�μ��=3�=5�><h�=y$<��k=�	�"��<���n��`(���Й=��w���Y, =���=��@>�5\>U@�>��,>]a�69t=���=��e=���=]�=zn�=���=߉u;/>Eb=t˕=d�����C 3��o(��	ѽvk��M�z����=�F9=UW���l��G����;$��<[߽(=u80���_�;,9�F'~�ڙ���=C<?m�<E�&�!!�=8f�i��=4��;b�|>Y�[>�1R>�R.>�ߌ��qM������L��`�;#9��j��O7�[:���<ҕ������Z~����g�ʻ[� �nʄ=�1�==��@�A>��ؽ5,��H⽻bk=O,���l=�H����>_��G���7N=6��=��L�p՟<Z��=��>����@�=?#�=Iҫ=I��1��=.(>��<�;��`�������4���𼭩�=��t>L|={�@�k�<`k�=�]�=�7��2(�=�O�<�5�<�zU���(�A$׽�CŽkd�;�$���9>������=�5�=���=p,Ͻ���=C��<�]B=�L���Ҋ�a�*�Hp��ma�6�*>e��=�:�=̶J>�9n>~ڃ>�q�=��s>���>�)->I�=R)>k�='�=��=k|���>�>[�t>RԽ��=h��=�'>Ѩ �r5=}�A>XV�<��X�˼ٽ�����<R���½���}V��a��j�=8�<�����-=E��=u��;�c~<��ýZ�<�m,��b��^��	����A����=&?����A�=��<g╽!���?�=�b�=.�a��4};G���x����q�<ݾU=�G��:�U��	=�����:͘�J��=���5 f��U��t4i>��=��c=��=w���c5=u�=���W�<��=>�b�<U80��>�bI=�Y�=E�����<?�콰[���;�r���g������j��P�=�?>n�">#���D�B<3� =�!>j�=���=Ã<�٨=����@v���<�eǼm�>������=���=�<>�DT�^��=S=t�=�
A�x�K�}e�=��=���>�Z�=�!E>��>7�=e��)�<�-�=��x=5p=�L�z�=�>���<���=���=w2�K�>T�=�rQ>�0��^2=_v=>�L���fl���=��<��:���P<��ȽMX�(F�vЖ=��=l>kƽ�p�=�k=�B	�;��Tͯ<I��=�"B�<���΢��(�f�	����=�W> ���/�{�/=��*����Ȓf<�_=�
�����=�'>=M*>� >Z'>`>a>J��=�A�<��;�uɼ�Rz=��!�+%�����<ǐ�<��=e�@=�R�=���>��>��>L�z>��=��3>)>=�ƽ-�=w�<<V�=��9���=N��g�w�;��ϻ�k�X��?�'y ��� ��;���;����ؼy���d=� >��w=�ϐ����=��>�<�=�������=�>�o�<��8=��=�:�S�Ž'��<�!㽤������묈=�P�~�|8��J>c�>�<>e�2>Q�>�-�=�u>�gy=�a�=/����3t�׽{D =�q9�N�Ƚ�n+�0�=|�x�\���4�����O1���d��1��M}+�6]�S`A;77L���4=�؇��R��ӣd���ٽhe	��4���(�G$�k�7�W�ͽjƈ��P�;V�5<pÕ�P�3��u�=ߏ<;~�<h���;_;kY��8*O�����m1����i�ν��X�l�:|4=�v�=�p��/$=8Q�<�|<R�*����^��=��N��{>{tC>5�)> ��>re>��p�Y�z=��7<�>�K=u���l����TA>��J=o2��0�<����/�}�q�3ꦾ8A=�ٽ����A��=i9�����XH`�̡Q>�]��Y�=@�ػq[�Ky�ե��)Q5�!���f�)��"�i�2�������G=���(���8?¢�oP<�d�=|��=\�?��>1rv�8�>�_l=�S��A3���|�=�X�>��	�"ZվM�ľ�L۾{Ğ����B0=����>���F�=g��>m1�w������>+;���(��d�;?�]	?#��>��?"��>Iط=|Ѻ>JM�>�վ:+�<�L>u$�=��ݾE �> ��<������Ͼa/���ʽu9Ͼ����1���ܾ{���'��	]�%L�E�?��>@�Ƚ">wj�>��>dp]>���>@�.=��C���>!5�>��;�>�l>� ���6��m=�6$�=�Y����G��=�>;2t�!��=�i>H��ާ���g@��,��B��=�B>��=��Ҿ��8?�s*�*z5�b�_>�?��?��?'
�>��&�L�?�����z?���Tr�;��i�>�r=�h�.�����K�1>�/�|�!�����S��p�?y4�=om�>��	>wrQ>#Cپ���s4��k=��n������<��=2���G���d<��aD�v:��t�f+3���¾�q=A���64������Ř>�w�=�$=���e?u������="�>:x���W>d5g>	YP��83��9?��>,��>�����<�ĥ>�4�<�7>��t=�	���'���f#�����_���<��x>��\>B}�>ϼ�q=�_>�｢xQ>����-�%��i�>8��F�)?#=�>��=��"���>�ĸ>����>{Ɔ>��=_�Ͼ�K���-��8a��l�Ǿ�2��O>(�H>L7�\� >���>�B�>�8�=���� ?��w>��@=�P>��v>\�\<�����>�[?t>��$>���>S�<�zu���Ծ��_>a�CX��v/��؈>�eþ#��7�!��Ӿ����B&���8?֘�=lV����=k�?�7�>z�>?9�> V����>���>�`?{�C>�F?O�=�o�>#���A����L����>!��=ٴ�&��=bU>'�?>|.?>5�8���>7fT>f��>m�]?O6'?0�����?�;ʽr0^=&��1��>�p?�w�>޶�����Qq���jK�R.���-���l����&ľ�FX�8�>w;>@ޫ�m�<����>���=
>�w?o>�qɼ�U?.?D$
?l� ��%(��j��* �3 ���R?��=$���F���nw���$!�=�4��(�(S����>W�?
�>���W�>8�3�o�<P��>���� �M?���>��s�	��H~����ܽ(�<=[��ECO��b�>Δ�<�쀾�4h��C>.;r�6=�f#&��:=t�=��%��H>JK�>rw<���>/��>���>;�R�/���e�c�5}9=�4/=�0����ҾF�;�Ҿ�������S�۾S��>ڹ;SN >V�A>�x=��I��'^��qǽ��Y�eŚ��L��/>x>4�}=�=i�>�֔������*R�_qþ���=tH�m5Ӿ�1?�M��K���g�[=r[�>!�>י�>�Ț>�-T����퐾��B��hپ��V=�[ּ wϾ���>��6�����K���>	�?Ν�>�H�>��>�%>�:�<G�>l�=����5���(�ԙ�=;w��+�>�msF=�c�>Ї�>~��>��>A-׽��>=���M��jͱ���O����	���n�=q��=��C�n��Aֲ�h/��N&ľ?F�g��e#�u2�ݜs��Gf��߽�>nt�KD�>mh�n(ľ�i�UVK���u��2�=��žB	�=�r�>}A>�ok<˄|>J�:�ɩ�fà>g�.�F?4��>U9K�m*,��BT����9��6�>���>��?IR>
i�>��<���>���>ھ�H�?�>9���;d�����gO�;.Q����>��!>��K�Ls.>$��=�Ǔ�)����(��J>	5�4a��۱ὧ�M>�G>M�T>,j=��>v�Z>/�=�>�ZT>X��������k�tݖ>���������Ѫ�>9s8>A�>�֌>�΄=?|�ᦦ�sc|=��=�����[�2>�\�^ C��=+=L��>�F?=��>�`�>�>�L>S��>�>�΂>[�>i�9�5ӻXs	?�R��>?�n�>������� 뾔���+ڻ����>�=?���>��"?A"�>U�=B�>A�>�ԭ>���X���A?��;� b;?*b�>pr>Z�|��]�kT���c���1==n�?j�=fT=p��>�����<q��>w@�>D�>���>�e(?���1��ܠ
��4���@w�H���%>����n�>y���v���ǾOm2��ž� D=��n���_�]?Žo��L�?x��>��'��<jv�>˵�>�>�a���>5os��i��Q�>��2?����u4~>W��>T�>�.����>`o�<>Μ>�;.�K��N�;?���>>����нNM�M��=O=�m8?�M�>%	�>���>�Ә�L{>��?ȏ���)1?��3?��׼�ӥ�+�H�����ھIiH>Q�>�m�>��!��u��)��8&?R*Ǿ;0$?�ՙ>'s׼��˾�T\�����8��
.�>���>�'?Dӑ>�a*?�5??m�?w�?�6q?��>E)?���>ӄ>Ag>��?;�?��z�$}�>���>5�?��ٺ�>͹���>iJ�>�F���Fm?� �>Yʾ\">��=񁛽:�1�W���`$ľ�o���ƾP7�<B�>54�=��$���>g�3�,���u����P(m�Ϫ���h}>��A?_uF>}JQ?�>�>��u=��>���>B>�G���	���-?x*A���>��k>�9����=�������d����O��>2�U<l�b�w?	P���%���s>H��>M�==��>&��>>�>|"?4�
?�Ԗ�T�;���[>�Ԙ>up�����>��>0��=�@��0xC�mĥ�됱�U�Ծ�[̽rKv�ϢK>�f��#h,��4>�������9��e�J-�<eݐ=�ܽ��=!��<s)\���,=��
=�O_?�b�>E�J�}��>�b�>�)?�������>���>n��:�>ʾ�9����>B�/=��ݼ@0�UP9�:���[_�D�����k �%S\��`�=�h�<$����#?��)��@����=䠠���>��>�*�>AEz�֚�>�����*߽a��Qn��TSW?���>3��\��sG˾!�/�-�̾�U�=�&�>�_>Kɸ���>�ھc �:�>�վT�j?�E�>j�̾�߳����<f��3J?C�{<L?Mx>���=��\>���l��=��þi�=l���p�=� �:>�y�x=�-�<���A>�pV߽�A�>���>��,=:��=�n�>�<�-���9j>�\�>��j>Y�>��>U��>R�,?��3?�&?���x	��3h0���?z`����?�Q?Mz�=64z�Rm��Ҿ����N����վC�(�������P��R�>�[?�?\�T=�_?4�%?�<�=a�i�=|h�>�i9>�E���\��H7���5���Gd��~>ʆ$<�龖�?�3��h�ش�=B�>ڣ?f��>�~�>'�?�}�>+�>���>��>��3�����7��a�<wм�;���O¾��ɽ6�����}�H�����>��j����>e����{�J�>l�=�����"�>�fG>�Ū<�h�&2�9	|�������;�����;Ц�����=�	�Ր2>��`>�>0�Fԕ>i*�=ԣ<�3t�S�<�P�<5w���jc���p���4>�\=��b�q��=��3?s`�>V,��mN=F�>@Q�=����1��=��>����?�m?��>s	�>�q�>:��=!q�Z'��m�k>�}�J�¾�W���ӽ�¾Ɲ>=�{>
����5vF��?6�\j�=^�����������u>��9�iT"��ҾX;�>��>���w|�]�/?'t�az?��dN���j�������=�cо���	.<��=5Ԝ?�ɬ���\�G���(���4?+�V>��?v,�>���(섾�ɥ?��U�k��>�(�����q�v�����ݢ�S�=vY:�֛4�x ڽ�k�>���E7�==,=��쯽G����ɻ�#�!
��<�p>_��>Qh@?x����@��?��_�&�@I%H?�z>H��@�>Oq�U�пS��S�1�&�����W���ܠ����%B'���Ŀ����>g�?A����唿��>��?��?��Z��+?)ߢ=#N(?Rc$�C��<�!]?o)c?���٠�P&>�;m_=�=��H,N��l�<:����o>�F���~?�8��$�'���8�>���?&|��8,�p�>��>N��L�?IR�?�gU?�q�?Sʆ?��k?�Ӿ�?��վ˒����R�� ����C>�Z�(��Vq4�b�?�b�;�����>'62��@i?@a�>đ"�))���𾽎C��C|�
ߢ��J?u�>) ?��4�B����>��?���>v��=`�?��? �`?*j�<��y�o�.����4?��w?H�<��3��D>L��=��<�Ō=EP�?�����NC��9=�҄��ɣ?�+�?�7辸�ݾ���<w�q?��ɼ�f)��f?ՙ����?��o�3�%�q�?�W���|ȹ��V?����i�>3V]>�d��_�>x�m>��߾ͥ3?()�>�}N> ���@���Zv�?�dF?4W>q��>�J�=�5o>ŕ�L�Q>t�g����?��8?�`�%f!�Q,�>�����?���?�B>�'��G���8?��Ͼ�DX���w݀?�]>���'�O?��j?	W�?Fk�>�F9�@�t�a�='�"<�ʉ����?b�>�S�E?_I�=`�����ؿ��D�
D>0�)�N��>L� ?`9�%ɑ?�s��j�>1%�>��m��g�>��:>E����S����1?+چ?Ι�GE?y �KU�?�y��;D?��F?�Ľ&F?���>����8�>��5�۰s���$@s���/��̫>=�b=n�B<|ő>���wA%@�?>�9?9��<]ٳ?����w����t�u��?�3�?SJ���|���>��8�v�¿����7?�$��S/?�$i��Y*?����*N�H1?^Cn�w�t>fa�qx�>���>C�-?�pw?�� >6}����+?�=?6?���g�5����I>گ۾���ZQ������H�vg���=�>��k?)����Xa?�勾i�a?�،?~�V��>�*8?�T�ϕ@X�t��S�����O�=���>�^���۾�U?x����.پ���>V¬>p��>Du��X���>+�?%�`���?���>)��?J�?q�?��l?F��?�%S����=/�ྂ�?*�9?�����4��R�����h<���<��@?�f��?5��>���>�ο��P?���?��E������>S����?��1���n�D�?�)[?p�6�@��1�־���?˦�?}5r�4�J��9�<P�ֿm5�?C6\?#ٚ��Z�[v���[>W��?'3�qhF?��>�Im���>����k?}�7�a1�>oW��s�C��d����y<�o�ܓ#> @��P#нmlS�".?y��>Šy��U>�է=GX��q���-��o���f�?P>(߁?- �>�2�>b�S�����V���{�����>���=��ɿ��=�)�=d�>����2��=��h���?���������������6��H2v�c���!?4��>M�,@#{޾J�B��>T�?��㻛ލ?i�\?�O��!/?|?���>Az�>�m:�ٖ>����r;�i&�?ym����N?>h������F���V^����?�̂���>��?뵓�(�@;n�>tX0���3?�ֿ�&���x�?�
�>���?n�)�������h��W��G%? ���՛�$�V>ok���n���f��*����zv��!>�x+����a�*>�s.?�f>ʠ��v ?���=�7Ѿ}pO���L?`>�=�c\=�����w���?�Ԛ��k��~N�?E�?�Q�D�?WdA>��?�V��>f�?� ?�(?��ҿ~%��B�������>ǪU>�P��!��>e�{?�3�?Y��?�U6?�_�>Ʌ�>�� ?���?1j;t�#���_�z�M��x��.����]���?5G��.��>�U��������?���?7h�?j�?��>�44?�`"?�rJ���=W=I���2�V>���w�>�ƾW�O?]��=��>���>W?�_?�?�.��
r$??��?;aݾ)!I?�B���tV���C?)�.���<���=1W?�_���P�O_7�/	�����yl�?&��>qǞ?���>�VA�W�P?C³�7�t>Fwľ-�\�@�d�W+�?`����/F�3�?" ??����?=+?�*�?[#�?�Wd?>�>R��?�P�UO�=ăf?d�2>L
X?YR)?n����B>��ƾ�:T?��?���16�8��=U����>�,o��j����@��=3oj?��?���?�?L��p�a�idd��`꾹!��J�<g��>x(��k1?f��>�=�?�������>��?�w��{Lƾ�"��b��� ����>����� �(1����?�L>䉓>�>&�@�6?3ْ?ȁ�>�Ee?��O? ���}>�>M�Ku�>I�r?u�?ߒ>>H3Ѿk�>��?p��>����Yo4>�?��4�Z����F�>ۿݽ{Y=*�۽x�-�儷�I�����>��>>h�����>T�?rH[>�	������EH�<�������@�<�=�MN����=���>b%??�q���f���'�у?l�?�P?�ѻ>{�E?���C*��,>I澾�K��k�bc���bN�� =��p3�Z�ȿ�>n�>֢u?���?' �>�%e���P?C�*<���	�P���q=K3@>�4�?����<`{?j�>p�8?�վ� ��	̾O��>Wr�:���P��ĿӏP��j������ې=i���r	?,��?)뾾��=�⹾�V��	��M���Ү���B>���?-�G�m!��6yI?]U�?=�$�bݾ�-ھ��@~I?�	���>�G�??u��S��?Ӂ}?n��?~?X����������G�@��?�m�n(ƿ�e\>t����`�����ф�.L�>
�������W?��/���j���?Z�M�z(?�0�3���u��Ⱥ�ԏ�59?�G�=l~���?#��(�	@�����k�RG�Ρ�%I侊�j?���%tK��뿿�^�%�p>�xY�9ڻ?�8��~�?�iY=�}��R�Ҿ�P[?�?��t%>oCҿ8��?#���ך?��2�ɩ׽��"'G@�@�>D+^�������ӿU�2?��=�?3�b�I�����G>?��>kjͿ.�g�T�2�x�ھ�\�=��!?��>��J=G�@�?��X�
?�
����?�k�>��=��a�k?���k\v>��t�3����?=��L���}=򑕽�)?:��>�ɣ���|?(@?v��?E������[�??�Mv? A >�h�����_�N>T_?uЄ??�>+����A��M��;��&���=��<Z@�?j��.Zt?�G8�u���@?�w��V���W����d�5�@?��?�yn?�>S�O�$){��t�Rڿ����a>�`v=Nm?T�=���� 9�)נ��n�?m/���,@��?խ�W�.���<�p|�?�����H>G�4���X�Ŧ5�h�@��Ay?|��>12M��C?s��?C-�>ͨ�?�?�Q꾳F�?2���:D?��v��y��*�����MI��"�,?��>�p'�����6/�?S�8�i�?�����U���b������&�
���T�?
��?% 5>I�?Y����y�>��>�=>���#Wv�J��>G^�!�
?��%=;?��8�
=���2k>�
>����=+�U���;KB?GHM��&��!�a=\%
@�!�?+��qv�>_`1>e�=7>ʾi�>4��>x �;J%>򒀿�Oξ/�o>��>mT��?J�n?��G���?�$ ?Є�<�Ni>�oG?fU�>�!�??���5>|���C�H��F?>��u�r��>�<��kp����>��?�o���:?+<��Zξ-�_?�9^?�h�=N�M>���{�>�m6��7S?�2?��?�Ž�$w>k��?�����<?X�ž�LT?#y��5<�l�?0����-�>b��;�J=�	�]��>��	��Ȩ���d��nC�x����7>�ħ��>�=Q=`-��U�=�� ?�����2?�؊?�f��]?ic;?N�$?3�t?h?�>]Z��<A���<�2�>6�:>��}<g��>6??>�>߽�Ƥ= ����^q���=�F��0�a���7�}K���>A>>��S>(>I�?W��>T�>B{?4G�>�ș�S��\4�>������wҾ��">���C]��^R���>����.����nm����U��>��[?ԮN?l�?z��;}`��r�n%w��	�>������>(�ǾD�Q>���վ�	?�1�_���&��(�<>� �>F�/?!ދ=L�O���9��k��՜>x=^>��+?�5(?�+�>�Zf?  �=�{��J����"D=�lp¾��?���>6� ?���>a/=ݪ>��վx�	�؞?`���U���������<���:����i?�_$?�4��q�=o?l̆��/r?F�����[?d(>GWJ�L6���Ӿ(�v?�k�J�&�>G�&�c���P�¾���>���>�T���>"*�<L�]�9�����h���� ������9>{�Z>�n�?ۛ$>W0���F>��< �e�c�Q>�D_?�H�>�������>�Z>\�=Y�O>6o>Ҁ�>�X�=�1���n��WZ?�V? �U��1���@>nT{��.`��U=�^��/;O��H߽ٹϼ=��=��L
?:�A���=�dWh���>׷�>�mc>�?�uľ��3?��c>�s=?d	?��ƽ�
?_9�>�>UG,�K�ѾS@��-s�����&|?���M=pF����B�=_b��a[<�O�>>?aQ+?�u��R\��ŕ	?�򊽛;�=�*t?��Q�`�d���$����s�,l�\$����d��>yw]=6��j7��W�>��>�����?㗱=x��>m�=I݈?<]����>}Ez>,;=�������=�	�g�h��k�P���4���=D�Ͻ".�.}>���坾�֎>�y?z�n��׏�
E;N�����>(E>�S>a��>��=#�=>���cͽ��}�h������
�⾕u��C>w�����p5��"#?�.�`�/>�ꤽk�O>��s=ʀ"?�z�>�9����m=�u����>�����>���_�i���Ⱦ}z$�x���I�> Y�>�������=��=Kw�?k�=��C�dز>��F��|�>�D�� ?�J�>�b޻e{�={�ܼ����=��"��r>S\"����1�<>/s>�E,>�w?�q�>�S2?�?�>����+|>R�>��>�n?��� 1?OO5�ʯ׾�1�>^�g>z��>nf�>r�ӾZ�o=��>h��=��?,��>2�����o�-��5FS=�W޾/� �ui1>�e��M�Ҽ��> n�>#'�>T�?^��>�Vk>�&�<wBܾ.�h�/�>�f�>T�(?�we?�-S>�}	�Vİ���>|��>ޱ$?����A��׾����Ȟ$�^���-��R.پ�D]�Gg�����O����P?�g>��K�nV��@��?��>x��>���3�Ⱦ�I|?�[.?`�?�#??�'e=8�S>F���5f�>�6�&ű;�/��I�>5/�;C��)ٽ=�(�A?8�<�>}�G?�d���L0>�޽��о\16�G,B��` ��s,=���ѦW?ä>���>���><pw?F�>[<�?wG=�=8?y+ܼ؂�=�&r��JA?0��=�[?�����P�>�#�=V��>��V>~��=5G�=�����AE��|��w�>�d�$�>��?-<>eq�>�{�>�g��GQ?C+�����>O�Q��?�8��>�s:9�W��i�i����f?v
�����>�:�>�W�?�Q|=,A�=������T>�oϾ�� ?h8?2���6���u�=3(����=ygg����N���Q��=:��>�V�>mk������H���J���bUm?�����^I?��?��Z�]kz>|�%A��:�>���T�`㐽�L���?վP�d�ssξ�
v>ɤ!>Oݞ>'����>�p>s�Z�p?�m?�6���7���&`��� �B�<j1����x���
�"�h��-�L>4dL��+6;a^�>2>���>���l�t�XW�>�$�Sbۼ�#?�U��˅?����{�C����=Y3?�7�;��1?4�Ⱦ�<�&�>R*�=� ?��̽)�;�:�:~?>�??;����>�n>�p�f�-����r�=ꄛ=)QR=(�R<�oU��T�>ɟ�>*&?��[?m j>Cw�>�T�=�?�v�W.�B�����=��/u���¾cD־?�i?���7&?�K�=iY��a����=i7�=�r]>�q��ں�>^��W?��^� >��P?�>�S�>^9?GA\?	!$?��A?I4�>	�L>�&"?��=h��>�3�>Ae?�0?y�}�P��U>���ܾ�Ҿ��T�l��>I
.>�4�E�7>@��>>$�4�+�ʛ,?���>�I-����3���H��,�������F>C��>� �=��9k(>>�o>W�-�/J{<���<y9½�V��ޖ=���>vgY?��BI�>��޾�j���W?���=��(�c���=վQ�<�5�嬦��kF�7\K��~<�|>�P>��p��uH���k�TXQ�9��z8�-V�<���h c����>rA;>y#.���T��H�=u�?�D^>�?�&>�մ��4½ٽ>�h��>]*�<쵾D�E�Ts+�Jx��/S>=��?ʌ�=<?�=<ؾa^U��h��Y�?"{��Ũ0?B�K�i�>����'��`�>I�0�(����TO�ڀ��==w/>����La���Y��}>3���c����c	?D8y>���H+��>������=��=��L��y>�R�>�$k># �>tte�"8�><E�6ʁ�Q��>�_T>>B>*�R?��9�2��=絫��>�>�/��%= ��g��}�b?P��=ĺ�u.����	��ڸ��N|��)N�����a�=Ëy�mIܽ�/=�����5��~�>~�>�f�>Ӽo���>,kv>����M����>r:ӽ�o�>���<�6��i
��?��K?c1>�v>Dn$��c>�n���H������Q�Z>AA-�̚�?�TR?��.�[}e?��E��ڊ=�Ԏ��n���/��>	gD?ߵc?B�=m��*@�=�_��[�?HǤ>o��=�+b���{?��B�?o�)?�n���=�<q�=$��>��>,?�� ���d>�`���RN��m徽Gn��/�IH��e�>WN�>�[0?�^�=1r�X#�=	��>Ec��+��=>֏(��y�<��F��>;ˤ��L�M��˶�=̲&?��>bE���D�>���>�Yn<J�]>w0i>y%�>�8=?`�,?1e7?�Z?f\6?���' ��5j���>(j�>��=>A9��o̾�ٮ�>{�W,>�_�=1H�+�����U�J��=s��>�4�=cF�>�q�=1�K��e2>����$>��𼜎���G#��+�����j��� ��𿾶��=8I�>�*N>,̍��#=�D>�S	�V�ʾv	���5>T�P�aR���d�>���>$�?@�n>H	T�nG3?վ�<�m�>�!#��G�>�>)K>z�Ⱦ�˱=��u>��?ފ.?�0?��e?��O?��-?E�*=>a}>��=�HO?7'?	��<x�>>\ >nf�p>va7���̽o0���w��M3�=jJh�j� _�ݛ�>~��h}��a�	�d��=��¾��>cm���`L?~aܽ���-"1��>^��̵�?j'�?چ�6�#?�א�)�t��`?�C�FN�>;N+�6�?Dx�>�1?�E?�����-H>#�Y?�Zv>6�>�J���]��ї� ��)�>M���'��&>Ц����]?�6?P@���@��א?毓�Is�>��>6�g?�m�?��>
o?�z>���=*����Z��X��T��+f�=��?+�j�ʎ���t�����N��ߜ7���q>r�=4x;�1b�sEX��\�^졾yܪ�����L�P>��C@���u�R>^2���9�=XG��¾�=?J0@�>��D>��m�l��>�;�����a�������=-���-�߽��>$	L?#E�����a2C?uiϾ��a>�j�<����슰<�P�ۮ��d���=M5��Y8�/ǩ���?6{d?�5	?h?�?@-�����d+[>L�?Mm2��D����>闶?O����S>{�򾗩>N�\��,�<Ᲊ���C>WӞ?t��>ЧO=�� ?#�8�F�ۿ?.𿸸�=�Ĥ��/>�b�?r29�*.N?���>�z	����>��?�Ͻ����/썽6�|>�����m�?��?�%?HH.?�5��"���q$?�o�>��?���>|�<��A>G!k=��:�]�>�Cν���Eo��Hz����O?��>al*�55>n�]��#z<�L>_��=��>��A���=��!�{�]�[�7���?wh�����=����`%�;�2�c|�	~�?δ8?z U>�-@������쿍q�>F��?��	@KJ�G9�?��>) Z?n{ܾ�~�-|��K��̣r�Vt�>��i���=��=̯?���[�?�PX?P�?�;Z>�m��㖿e\�=��A�iЀ?��Y?9�"?d�T?RM�>�<?�J�>s����f�m2���>�����:��=���=Rʜ>�_���ʾz�(Kh>�@�����ӻ�?2�q>a��:^�=��?M��νܿ
���Us�?���0� ?�
4?t��?�܈?�??�.�?/2���>Z�;�C��]Z�?>��]C�?B}�??�Q<��"?���<~�t�+?9P��T?�9J�B�?vBn��z�>*�?J��?�� ?^�>��#?P���H���[�MJ4>�>=�֢��7�L��t��u��>m��:B�p>� s�1�?�.��{�=s?\܏>�;-���>k�J?9��?O?@j����k?շ�� ��P�?'7>�[�"�?9��=J��>W4������j��Z�ۼ>�	�jz����>m-��ER{�B7ྛ��&��`?H�>�W?!�4>!�Y��A��+�:�)K�J̾n�>�-��g>S��?�y�=�^���=��d�?����Xv�p�&>���>Y�����=�\Z>��?�ǔ?*g?Dz�?!p�?ȶN?�Q}�-^8�7C�>��?l�>=�
*�,���}y��)��@@��Q^?�NC���?�4�>��?������=1�����|=ى>�|`?�G���>đ�?�8=Iս���%?�k�~�+�@bt?&�$��G��GU�>�q=��-οj,�i��H>qI�=ƺ�>��_?A5�Є����cT �GǊ?�K�?�,1���e? �Ǉk���(��=Zo5?Э�>�;�>ҡr>�5>��S?a�������Q[=Q�>ť��D���6l�*�⾼s�>z�½e���*��b�?S!?��>q�$?jO�>�ba���|>�G#@�~�/Sq���	�a�e���T?v�T>�AK> .Ӿ=L5��_��2:������(����&���y�x�d? ��6F?�彐��>�显ޡ��]�<�I-��P�t>�V?#���<?[Z\>�D6�
V>!ƾ��x�M��?|kM?��%�oOc>b�Ͻ�yZ�zO]�/~��ё��ѭ���?�j�?`���9+>��>�=�
�%?݁��C�j?�y��|u��0Q�n���+�>2�?](���怾ebT��c�����{�F>������.�P�ۅ=?�[��8��`�>�,y?�Ĵ=����>T�?���BhF>���>Af�>�h.�����W�u*?T�t�+j��GQ���8?gd?��;�Cr�>5�6���?AM?Fo?�|@?�#���ҿh�>?�H���@�����?Y��>�*>Z�?�t?j�E?L�A?�2��)�4?�ݾ� �|0?Z�-?��v?�>�����i<��$�IR��!�Oڇ�ҁ_�E���?oP>e>����=^I�����G���\��Y@�U�>�;�-��>ߖ\�<�~>@G?��=��/?���N�E?�����f俅M{�8��?+��}��>��<��?6'P?#�g?{��?�#�a�=x����*�^�&'�� �R����=P[��.�¾ڏ2>X�6���⽱C����!�;�Wp>�^�;�˾�L�?��^����� z�>�6?��ؾ0�����ھ�b�?1��T�>��=���?N��<��*?	P��L�<>|��=N����=ǈG@�>/H��N�=�L>�ғ>��/�Nu�����>/ϣ>� ����d�>O����!B>���?B�H?.!��bo�Zʈ=8���z���۾I�Z��������>;����b�u�G��C@��=?o�:�+k�?����B6��K�
�ھ�r���$���?�h�G>��9� uF> �^�B�>?@��?N�[?���>��?B�~>��?
�>��?>�<�?%�j?��6?�՜�v��>������C>@��m�B��_1����?m�D����d�?(��>�	��2���8��=�ԣ�ΰ�c!z<z.���r��<F��>L�k?��=��p���9?��=^�`{�PK>��>��Ӿ������?ƀ�أ�SN�=kd?�þ�������Ƣ`�slO?�T�?fP���>�����R�v#�������>"��� ��>�S�;?���D�q�}��m9��E0��*?O0?͢q?浙?�5�>u���+���=�� �>ꣷ>@!@�^��ѧ?�<���>�i��D�y�?j�>��F��`&?o�?��>ٵ��z�[>��=� �>�嗾_b�>�?Y�&?��U�;J?�x�=�9�>�Qo��z��30�>���?>�\:�?;�I>���?_��Xk�� ��>��?���9�)��y�?w��b�Z?~��=�滿�@�)�>J4���?f}?&U�=�p!?�����f�g�?��?�?�n�_(���/j>��)>���������l���9f�?Y���2����>����b�����>�3���R����='?,� c�;��vc��
�	� 6 @N?������%�	�22���1�7f�\0;�$z���@=D�?v2m�K��H���cT����X��>��7%F���{>��Z��F���Uk���󽁵��kQ�x�>h}�Hh��q�!>0#0<��=�\�>E.�>n��gP���2�^;�>>c>�j�>��>����>�?����������@BG_?#��8��?�Ƀ>y��>e?���2>�a�<o�G�y!���wC���l����> ��=���>|)�?ڻy?�e�?�B=���>�|�>o�=i)�3��>G�v?�kb>W��z��&�?Vc?,B�=�?,
>��e��Y�=��q?u��>�ބ?2�?m`+>H{?M�A?u. ?%IĽ!~���,����C�:"�����T ��W��[!���`���?Dyi��0>�	����>Ǚ	>��? G
?<�߾�.h?{	��I���H?(��r[�>vC��)����`>���~���=Y?�a%�aҁ�����]kR?�
#�c�=�e �����Z���ϐ?#�V�3�
�r쯾�z���?(���~���z��ƽ�����?��C�B�?�KN��l?���E?�Ӿ�?E��>��?�?/qk?L�>5�>�H�>օJ�~�?����Nڌ> �����>=�?g�?�����܋>����ԍ ?^��9ۦ>���m>�?�\���>����2�{>�v����\�����?R�,?�蓽"
��/^>k���c�ü腜=i��:��D��W��I��L6��b��1��ki7�A�0<~���}Y���o��>�;�>đ?>��?���<Iiq>�Ǎ>
^>��ټ%�j�茥=���1��ܔվ�����7�q�ɾ���FqD���0�L������i³�q�n>�����L
����#��>�>.>F��>�C#>���N��=��<m���5B>BC->z�%>������>�KK>�6>j��;+���������ྒ�羣ڀ���>�I+�<�!���a�q"b=��>��нYg�>�o�>� �>P��D|�=q�o>��>\�A>�%>-��=.�>E��;އ!=��1�~��=B���'z9��	���s=8R�>�3=E�J<�*[=mE>�/_�����M��}I�=�p)�b)���/�l��_`[=}�%j��4c>��?>�r>�K�>�v���{�>l9>7�>�4�$��i��<���>%���K̪�g8�k��=�	f��Ҿ�򣾕����>�>�F<�y�>��r>�Ec>��x�:���^żd�9=3}|����h��p��={n������M�=1T�>�t>��`>$�>J"8>����}=6Da�oi��Ga��[�,�$��</2ٽ��.=�|[>=�=�Ў�|�%�<]i�+�Ͼ��X��J>�4����#��|/>(�N>ܞ>�-�#<F=U�!�Fc>H!���b����ʂ2�P�Y��|�������]�=�*x���=��>|<R_>�g�=e��=�=Q>�=�1>=+E>J*=���=�7=���=��y>�GĽ
=h�����>�O��>�R��0�͔���y=�/`>�ؽ��<��!>��L>�܅=�C0=�`w>�aa>�`�=VE*�����y=08o>���P�>���>�/�<�->f��>�A�>��; �O�9>s׽-誾�T{��M)>�$���Ƌ�	b��*->}E�=_3�=��>b1�Ų���<�t �>O2,�Hy��T�=�y��>�t�;l�2>�V=j��>S��)^>>N��%'4=���=��m��b����=�;M�O�x�p��r�Q>�aҽ��վ��C�A�<>(�>>��>���>��Z>I�ݾ�I>�y�>��>��ʾ`��>�k<0=�>��C�pԷ<�B�共�����(����x�y4��&6��D,��*Ӿ��^<4��i�2>��`>�n+>$|!��U�=��N>b�r>�J�>ʀ�<��>�ҁ�I�C>׸�>��>1É��]��W����-<�����e
��M� �v�㾗�>u�i��%?�3f>����l>���>��>$����_>0���>CG�����,�f��,�j>��_pG=li�>*KT��!~�F�7��f.>��������~A�H�/>rd>j��=�/�=m!�>�?E�>�?�U?��U>E���+��>N��>P��^c��"�}R>�;T�Gg>��C��fa�=sX߽l)!��oy<���=�H�����<{�1ݙ=��ռ�D,�U�a�g.>-#>ی	��JK>�Lw>��;����!��j�o�䃽D�"�ȱ�
jC�~d��D*̽�ǽ�k?���A>^O>U��>�f�><(�=��9�i>���7U�<.E	�A�¾&t=���C<޵���,�8-��C	N>��e>,`>���>L�����н>������=�{\�:������y��<�x<%{�UQo��`��Sm>�h>���>�K�>��8>:ķ=B<�^>"��@#>[z=ƺ��L����RF��sR��<��'��������Ǿ�b���\����i�����վ�I�>D���=�*�-W>����z]ټ�8�49�=�2><�j>������FV�>�>==��Q>q�9>(�>,N�>4D>�1<��<94
>N��=z�N�p�ý)����u�k%�=ae>9r>��>�>a��=L�>xJ>@��6>�P>L��=O�w�r����[��샭�l�">�\>���5�@>�6�=h�ü�+{��K�A�>[���+���z�u��Y�>i>�{j>'�=�>ۏڽY�&=�K�=��=6<5�@���F��e�=�����֮<��<x��>�> N>�qq>"�e�Bk���k!��T,�gU�<;[�?j	���>`b*=)!�;K����>&>8�>+��>�c�>8�T���>\(>t�>�##=�0/>��>Ms�>:��=;3"<�e�=wgU>P�'�K���M������ʖ�(����Jh=����M�G��9>�c>��$>��=�V�=$F�>�G>���==Ԕ= ʩ;u��>��I�ZSо�������g{�<e�2=No!�����;��:8Ys>��=�Ӽ���>j�>l�>0�>kp���g����ƾ�����7>�]�� ��X��q�=P��m剾:>�Ȭ=��>X}�=`j��ۢ>�s�܏>���>a��=7[���7�=C*�>��b����Z\���>)�ֻ8�>����� ?%_��Y��<�c&>L�;=-Î���>y@>z�'>X��Re���{=@5�hʬ���b�%љ�:=��}ȗ=���>7�r>�Z?��/=��>d��>"��>�E>v�<�2>?X�><Bo�Ǯz����=����NV>v����=Kш�z�>r�>G]�>m�S�e�=?6>��>�й��J�O����h��=]ھ��
>_�ν���>D��=�?�>>�86?q�>b��>�?�?[�>��>��?�( ?5��>�ͽ�
=?�	> ڂ��Uc>}�>��>�²�b�f>]t�=P�>��}��/�=LП���>���7�i�ҏx��Α���f��c=�d����ӽ�p;�ZB%>���=}F�3V��t��`h�XB���T���sx�Վ>��=�I���m>��r>�<�>���=�h>�9?f�>wQ>=̘�+�=�tM>�~.=�$澊�x�A��c�	�"�%��:޾u��}�H<��ͽ7+����O��N>?�$=�>�g�>><D=+�.>>�~%��.�>�ʳ>(f�>��3Z>��>O��>>þ6��=�t�ᚄ�֊��b� ��h�;�2 ��g����뽎X�=�Ľ�.����>V�>)C�=}�a����/��>����+a��΅m<���=D޾"�a�f�>RI�>@.��|[�=#�>�a�>E���B5���$Z�w�=< �>��>�A�>aRQ>�9�={?����;�&��_"��ܻG���6>��q�dнI�?>�d&>�P
�J/�=�!?9J>w0i�1��>EɃ>��>뗴��pQ>2�� Ԃ>����U�
�A��&���u�	Q����>F�=����-�> ށ>���>�늾Nk���ȫ=�d >�<�:���q�t�:S8�������<L�8��$O��Y��������0�m�u>.�>r�=7�>>ˀ|>�z�>��[>d��>@<�TM��Y��j,������S�)���h�C��U�<w?7��_N>�a,>Փ�>�u�>]�>I��>`��=
� ?�޾O�>���>���>���4>=s�=���>�L�y����-,���~������,��/���K˽d铽��>Э,>�>�<w�R��>���>�y}>+֣��E�=c^�<�,=��=
���ޒ��f�-�n�;�׽~W���|~��>.����=)�<=��$�>Qpo>4�>�;�>��>�ñ>6@Y<tu>���>��>z�4�$J>�.��="�ν�@о��*��=�t��d�f�þ��->��<�I�>lZ��DK�=���>g\h>��i��=:�e���н-[���Q���.��Q�u諭T�y�(%�=�D�"@Y�n��^88>���9]�:�'=�:�=q�F>��/� >���`��u����ϽFP��Ծh(q��̦����� {��ŷ�=炭=��ྩ�c>a->��>��ؾu��<Xv6�ڹ�=���>Ϣ�>��=��W>�(�>�>J奺2ޟ�cZ>��R��c��X;����=w ߻�!�j3N��4��;�a���
�h�#?q����A�Q���"�>�����VӼұ����>��=le="f��M*�t���94>��KP?5
>F2��(�'�����}�=���G��%��+���]?7�+>���>J�;/�6?L��>��&?\]�>�t?Q<?@�b?�3?�>G_�@�<e�a��8*�L-�������ο��Ƚ�5E?�:��ق�2N����>��
�#�*? ��>�j$?��?^�?r'1?v��>A�>��>v��>�s�iJ�>��<>���>�揾Ǳ>8�W�୓�[�����U���@}۾��˾JlE��=�2���e�E��<߹?��>��6l@��Ô�B�P>$��?Z����!?�N�=p��>�?
��>v>�aR>�uC>�:�-b��{ύ>��@>���I���E����O=z׳� ��=N�=.[>�5��Sz������P�=���������a���c��E6?8(I?.�O?>�`?ž'?-?h��>ӄ�;���$ܣ>kB>�^���9�%��>� ��̶�D{*����=�o�XҾQ��O>ytB?v�ɾ��(?.
�>��D���׾`��<�O|�"�>�C ?W藿ֈ���sϾW������O�������پ�3�>�/��k��>��C>��Ŀ܃#>�h��+�>e���6�:��?ս�l	�/%>?�D:?�5ξl<5=�1=�o��Y ���%?[J�<�O�>���B\�>uɘ?�P���?�]>�h���m��>y@h>�����-�.�?�Ko>�$�eN?���e��:?9����f=�g�>�P�=���>�y�=���?t���(0��|�I<n+�=;a�>wK8=��>4����8��Њ�`,7�8� ��4�=��F�v�o�������E�V�ȼ2�?���>z����o??�=�i�>��>>�9�>�VW>o)W��T?0I�>;$?>�0�>N�?��a��i�=@��>j�)?��=y �>�귿�}�>����s��L ������<�a�����?�>0���/��?��?l��Gj���>Q���,?��e����?%�n?ۆ?�G>g��>a�?��>�>��#>������>�#G��S���>q��>��[>��_��2��ZxK>�>���^�>u؜�L�z?BwپC�">�2�ē�?l�;G�?�?k�A�f�J�����IG־\����\�־V���оv,���>Kҕ=�vཪ� �-��*��UΛ??.Ѿ}�>%�>��>2�	�=�\?u��=�;���>�N��c��>����a'?�⼘�F�
pʾII?����� �-���`�)Ę��<?���Ҳ�?R������>�_7�?�:a�<<�?��?(�<P%.�d)��SzM>Q~�=?&�>���<S�:�>�ʇ�*����3�R`�>�<쾓=�}&��h�>�W�=��,>r0>��>�͍?5��=��`=�k=>�2��ց:�f	���>!8��>�/��M�>�9�c�1��tɾ��<,�>R�+��>�E?O�C��Hʾ�i�Tƞ�� %=F$���Ī�>�>�<�>��=�����'8>�R�=��>�&���+�� �����!5	���4��h۾G(���B>޺�=q��>��>Z�	?��?�G��n#4?�c��F@�>1��>uA>��K��)�Ѩ}��>*��U�>�;�=��?oy�?�0?B�S?���>#���ꂾv��>��-�r�����"���Ⱦ��=d
���u�>̼�>���>��>�\>�~�(�>#�о?�x>��!���;>X��_��<�lx?�V)>U�>h'�=�!>.�>��=佾�aǾG���	�W>v����&=o�����>E�9���:���>�˾��8��dA��bE?f�?dY��>Gs>���?(�.>1�6?Ɠ*?�?�3?ᖸ>r+L>꾐�Q�'^����>�����E��Eμ����Gx?��O>ާm�⦐?	�?Ӝ�=Yh?�ȁ=��4�d x�Vc޾�7#������ ��>Kl,�����Jٽ��k>g�D�5�U=P�#��|�=j���L��5� �7��>��|�cњ<�ń;���>��޽���i>9�<������u/	�1
�=G	y���e��>�-�>�����Jّ=,s����W�L���`?��i<������~��r�>���8o?��(�_�u?Eێ>;��>�8�>a@�>�lF=�M����w?���>��v>���>���==���p�?�F>�9ɾ��O��=E�<�Q�	���/��8?Y�?/�нẺ?��
�K��>�U�?<�>Z�D>Jma<�2�=�:�>���>�c�>���*j��>�>$�;�#��
��o�1�����!���֓��F���$(���?*�>�Q�?�gt?:�ýJG���RI�{���h�?�7)����>�n�<ڟ��I�>e��0¾�>�p��e����h��ܾK4->:�ڿX��?��4o=�t���Ǎ?���k*��þny�=s�+�i�[?��j?�q�?�(b=��ؾE�6?�Ȍ?��?ӛ�>z��>�S?T�M=���>>]:?��<��@��P=���>9�>���>��㾧�X?�1��@?*3�>5?;��>%�6>֣_�*�*�{�t��$6���>�E�?��I�m[����?'z�=���>3I�_-?�}�>�8þ٧�>��	�����B�$��o�L�{L�" �f��>B!v>�#>[�>cԬ?�g?��W?[�>���>�GY?C�>�QW>3g?Tm�?��??��̽��̿D�>�B�>;�?xʅ�"�=RZ�> ?<=��/|+;�$?�;�p\�Ŷ�ߥ�-���k3���D���־�l�8�[>�;�s?+>Dk��f�����?���>AV�g��C!�>���=W��<�b?���>���kX?�ڽev޾Iݷ?%��=��o>��B��^3=��?�� ?�~>�# �V.���L�>S��>�.��#;>; ���þ������H.<
�
�%2�>�I+?���?�S�>�>�A?���>�?[m
>��t��M�>l��=�?z��>��i>6r����7�8pp����S!���6}�����)D��>��9!v?[����5��?���;8�7�?���>��2?�d����>ҁ@���^�3e��3�T��:�?80@?��~�@+��'�>!m�>s\�?JmL�"և=��i>��?��!�?�-?����͝P�z����J>q�~����=f9�>������ei:��?S���,��y����K�w�?�E?Z�����>X�>�F�?G#��˟�=3W5>��<���L.?��W>�2X��|,��>t�n?�D��;���z3�=��ɾ�z@�9ƾ�
M=`��wD?s��[?�B�>N��x8Z�38 �� �_f���3�UG
?��}?�?�=���	?T=��?a��>w$X>�L<�p���M>�>���>�Z>,>��>o�>����I�>ļ?i3��L?��>�����@�>�[9�]�?��"?T8?�F�?�.?)��=> Z?9��>�Bn��L?I(?D	�?@�U��ej?ǬL�8n(�������K�	�Ҿ~;�������N��@�>V�4��R7���?0*�>	䉽�"w?��=�t�=�	S?x��>o?��^?h�?�B?�_j��/��ߐ���!���ǡ�4����Kp�= o����@�$?	C�>MA?�V?'�9?�*?�� ?Dn�>�^?��<?*��=4�{�	k�>��=d�?�~Ž�X?D�d�TF�=�Z��T䖾�.	��Ož�hO?2����$>�g��#�>V�P?%�f��5�?�9�>[�o?��k���k�<�>�>޽�������P|=�*���`=�;��O?���>���P<?��%?ߏx>��=7 o>?�>U>N�1�Э�>��{>����y��	�������8>��B�tO�>y�E�$�R?Y #��>L>��/��<,>�q>�n�>QE?l?���=�����R�>m�? ��>�3��0p?�׹�/g�>�}7��ƞ>�З=v#M?sM��ޗ�~;�=�>D�-�&v=��n$���>K��52W��Q�=�7�>��<e�Ͼ�SX��?��ԏ?t��<�b�-RS?{L��K��z�w�L
���?������=w�A�|�L<�L���xG�7O{?�� ?���v���3i^?Uv�>�*�>`��=́�>%<w�E���B������䀿���boz�eN���N?gUY>��ھ.�e>�>��Q�=�H�Uxv���ͽ/��>�<�?z¾?��?F����>�&��NŬ��d�er�?�
?�뽾IML�v%@C9_?-S���Jh��P?Y�x�cF�h�>���}����ľ���<�i�k�Z>
`�>���RE�>�F�>ΦQ��֟>�\�?�2�>���=�jT>�v>��:>��?sM������O�>c]��k�T���g�VNV��W?�ق���I	X>Wo#������?��'>�<�>�j�>���<G���	�(>�*��o���_�>���?x��?��o?nE�?����"?X�=�QB��vb>q�=�` ?�9�����e��>p�D?��G�s$Ｗ}���߽���>K�?K����͚�F=1���lu�81����`�(���x�0?�����m�KF��YV载�?�(�=��?.��>5�˽j.�?��>dqq�$��>b�C�`?b4�$F�?�1�Z��>����iI>�����?A)���^�]����b�>$;v?�oɾ��>cc?|>��>�8�=ah?�t>��>EӐ���y���7���H���?&Ռ��8�[!n���s��
;lL>(_=lp[?ڧ�>w���?��YU>�(z?L }?ɡ�� ?�F?�����L��N���A?���Y�)?L �H=S?�ȼk�t>�P'���4�~h����l�R�
��?�bZ?�&��D��e�>�db>1ʾ�ԉ>ڎp?�r�=�Ҿ�c
�ּ?��?N���n�p��(�>���ʰ{>	9F�.�f�zj�<N�>�=-� G�=fx�=CI3��F@���쾀�h�{?!WT��I?ގF�K2f?\�>�<>p9���)?��??��+�լ�>�n?���bA?�	�>�5�;�{?:+���u*��[�u�$?z�i����>���>Y��?�9�>f+�>oa?��'��W�?� ?hp��&��Б�?�g�>�v�����0s�tJ�0�>��������,M�>��q>�΅��q濱�`�t6��ڜ� V�����=��>%@���$�>�@I?�����[�?�^����ǿ?տ���;��V>�Z�>��>mFN>�����Zþ���>Ie���	�������V���H̾�ҿ��=@\<_>��;���)��]?3_+?��*���~'�*t㾊�����="4?�>�?p�"�Z�A�g�2�m>3~K��U��0/u���'�H]ٽv�	��!��`>�z�>Z%���V�<�K?R�[?@��>�#;?�yC��򢿀����� �������ހN�<�������"�����4������>,��ר���ܾC�˽	އ��C�>	�=:vU>����>�B�Q1x?�@U��>����(��?�O�>���(؋?�IC�}��>(?�n�>p
?�����>���>�)?���>O;澞��>�@���]/�|#=�xT��"���?.��+�>{����)?���>ie�?s>1�Ū?�����>������L�h���6��%b>?G=�*��z���g�=��n��ɾ$\�*��>�:�>�`:?"ZW=�þ�5�?S��܄��Lj��?�*�?Z�����=E�l�B����c1��Ú�R�=}�f?_��<?�3H��-F>&���!3T��O�18h�)A�4p�����>�ȿgi�>�$*=��?V���?>B%?>��>�KԽr���)�>yr�T�3?��="tm�c?�=9��>*�����e�Y�ٿ#iӿ_꿅�;��p?�?�X��E?B��?���n����^=>��K���B�{��dF���F���F���W�8R��Kʾ��b>�RQ�V᭿Ա!�r��Ej>��^�ztо(�.�n�>����b�=K
v>�r�>������B � �׽"?��@wm�>� ���>��A�;�����Ն?��c���j=�;?�����b��WA���?����@��8�I���>r匾~F��h@����=���?��k?Y�<�H�>���?I�F?�Zx�<��S�?)�O��_�'F�u��]���+���
mI��>��8����d�����?�}�>d�C?S�`?4V�>� '>�$�Ov?:�?�|�>��>+?5o?a��>6	>��)��N=�Q'��P����GRY<o�y����X[���v?��ţ�0�1?Z>�qN>!&�?� d8�Jɝ���㿀|�>�e#�1$��XJ޾>�z?w�H?� �?�>޾���=k�:?�.c��}�K�����߾k�>;Z����\�?�t�c<?Y�l>�L�?�w��kF�>�(���?�5?�̾�r�>Ũ?��3��9E?��?`��<�r̾}��y҄?�o�?������?\e=�;�������c��e�>��>�!�����?��>�t�>̊?d&~>RJ3?�H_���"��ݾ�[^>3	G?�����߿�[.�bH�TZ?-��>#�0��C�>TN?R�?AW�?}`2���>on:���d=5�M>���%؇����>��-�F�?Ǐ�^�|��>�H�?��n??E/?'��=�:�?�U!?.�>=��^�(?�,"?�J<?&�>/-��D�>t7>Ҏ�W�C�����>���Z̼ˌ������>�0?R-��k��^������=�\(�G�b����1�#�>'�?��?�߂����pU?#}�>����t��$f��H �~����i?p�9���A?��?̈́"?�EG?Z)?,��?��?�nY?cDc�QH>�����2?�H�>��K>u�ƾ?�Z|>��?_@���7���?Eҋ?�ʕ>m�ݾ�A�>o?6W�?a�?��	?%��z�>+��?�̱����=)`ݾ@�k?���=!;>(x��70��1ݝ�$��(d��ܾ���9�?z�p?=$�>`Co>$��>�ih?�Vk?���?{8>�=�?vl�?mf?��M?	6�<N�����=�Ϳgb�?��N��
���׿l@�	�?]Ȁ����`d?��?�]�R!F�8f�>(�����*?���iC?I��=�헾���?\��>vv'����>tB���|i?�I���@?���u��>���ܠ>����/_?�!�?�Y]>���>�
?,v>N6y?����(r#���:?�g�k����=q�=�qK>Hn�l�� ��>��󾳴��a�@?X�>�'?�v�I��?�>���佰�!���FW����5�D�ۿ��ʾh�?�b?�[?��>��e��P�?F�>�AҾ.��<�?U�����?_>�3?��� ����@j��=��[�,-M�3��>-��>.`�<T�?�Rt?EZƾ=,�?(�k<��!�A��?���?��=,ʾ޼v���k?�*�>�h�?O
O��'��Aj?.��pQ�r#D��K��㏾���u'�<��}? 8u?�P?(�?�ތ?_�?j��?|E�?���?`�?"��?1?�"?�O<?�%�?6�Q>1)>,#�x1?�(��o��>�+�>|t�>pK>?�m`?��������>k+�?�u�>�6E>	]!���?p�?E��>)6�=�98>��=�}��7�>� ھR�>d��>��E>�mb�9��>$�.=��q>T���F�{?����]�?/`(�L��P�S>{@�+��|�P��i
=���>�ST�cTG�I��>��=(҃>�y.?��>�W�?�{D?�Z���
�>�j$�5��;a&�>�"����(�e>�>NO ���r>�No?�	I�Ӓ6?#3���=�o?)����g����?ֽ@�cſj-?f����>�|�?�<��s?<��>
h�*��>X�a�*ɔ?J� � ��>R�>@��=�R7?}[?Q��<($>�߷<�j�����F���??��>�H���q.���<��@շ���26�w���O?��<?>����0��ު=�����=��O=�,�^IQ�'�	�L<�< ������@��<dQ�=Jz�=zg<���˓=�Y�=>���=^B�=�=��=L+̻�U�<ӷ3=�z�=�=���-U��9�+Ag���1�H�&=X��;Dr�=r�f=*t����8=�>i�=��<�럼��1>T�6>��K>5�q>�1t>�pv=�~��t߭<���:B7=��=�F=����rd�=v�=�ӵ=�����/�F��ל�<l8�8�H�� ���yg�`3��Rt<�E>�J:>V��~M=Z�>�!>ޅ�� u�=i^�=2�*> w>$�:=j��=K��>(%�=��Q:L�����<_P<�\�Og��e8���=p�ػ�����=�[�Q�(��pҽ>J�}�׼+.�������C�D=tVڼ�<�R���'>p�>-9S>��>>zk�����aYV<��!�I�׽|	x��ȹ�0����3�<xǽ���\�콿�>���C�jg�pB>�>�G>��A>c
!< r��cKK�}�)�n�������*彧��F��;Ϙ�������=�1�=LX=�;>�ˎ=��=��[=��ɼ��=�\=6:2��=�m�="�>���=Gx>� �=�ǵ���	��ų��p�O3u=��>f�S<�'_��Ղ=Lޞ==F=�������Q�=!#�<�����������0�c[�a�߼
t=34����P��<�,�=�~�= ��Z�ҼA<e��=����=Y��<��t=��X���<��T=�b����q�g�=��=��>?��<����nb�'*!�w>8�P2g�ztټ7�w��?��p�=q��=!�E=�����*�=A��=E��=T����g=8�=	4j=�G����,>W�=\��=A.=>8k�=���<)��<�'�>��ż�"��T( ��>����g�B�/��NO=�"�=	#����>�7=$n=���=o��>Y�F� �=�{�=�5O>�/>��$>nþ=�ĉ>Nt">�k%>DAC>�E�>K�!��^=���;���=,��;��Z��+��=y
t=�a�=��X��>��=�m>o}�=/\(>j ��C�>ZTf=?:>p~����=�m=��>�ٴ�0$ƽl$���=5�����]�ܧL�|�z�x�X�D�ý��4�=�
8�ǕS�����B�=��5�0�?=�F���q>ȸ�=)�c=�G=�p=�� =��<=}j��d�ͽ.�h=��Ƽ�m�=�|��xn��O�;�%����`����1=�_=H�=��6��ck=�V�=aKb>di��Đ=��=S�=�0��=����Խ}��V<6�=y]J=Iy�>n �v���^�<��=����½R��Ϲ=/�=:�=p�=�&>(��=)�#>2��=�I>(��hh=�͕=��o=����SѼ<N����=aҽa@�O�������$�����f�T�b O=�������'��D^W�@+b�Z���O�Y^ɼ��=x��;�v<���=BB�<������{�p�ԼgAM�v��յl��M���=�S}��&��[�L�d�5>�S8>�_t>��>fN����?����t[�Ϡ"�8���,���1z�<�d�=޾��c�c��K��!L$>	�(>��T>�1�>-4�;�]�;�=|��=�
�=�����b��=J�<\��������<Xj=>N�=�8>��>���<�0 ����=��7=�=Yi�<1�ѻ�B��Y_�<Q6}=WV=�Ct���f�Y�8��D�{�r��g	�X���?���
�}Y>xW�h��k�D�
�N��<��g=�F ��A5=�<'�<�7��􀽣a��l׆<H;�����5Ƽ	�\=��V�e��};-O~;��<�w7��x'�n�n������Zp�g�;�㠼ȸ��gr����~�<�����Q��;�}���O�wTl�.q=�L���t�\z2>M�<���;V�=���=^���H������n=O1|��ڳ�U�=d�B>�,�=���=���=A�=����^'�;�(�&�a=�ڽ!ˣ�?Z1�⡣=v���}�Ƽѽ"b�=7t�;��<[�=�m|�E|�;~S+�CK���`����1<���v=�ډ��~��^3M���=�
>a�>��b>�
>Č`:}��<6�='e=��P=E��<�S�=�'E=�-��p:�<YQ�<��h=�3�[� �1#��46��w��g=z�����v�d¥���<�*�=M+�� 3��Ʉ=���=��
�gcj��"߻�g���9���&=��ϻ�=qk��=|�;�(�;�I =���=x�=6F�<�`_=;Kc>�;>`#~>%z�>�G��{;�%s��ٽ��H�k������cW(������y����ʼVM�tX��x[��p���)	�On��5�r=1\�<�/�=mDn���Q��8;��=�����t˽iE=|�
=���<���� 6�.��==@�u�0RμM=-��������D=���"�<�(;h��=m�L��}��y�9�Lk���q�<��ۻ���=X�x=��h=)=y#�=��<̏k�,0 =S=!4�X0���ҽ��7�`�V��s=��=��=:���8=��=5��<��t�h�O=E��=X>�ڻ��i<������4�սM9�=���=��3>S��=* ~>�"\>C��=�L>�>+Q>�Y>�/>�wO>}?K>Q e>��>�7)��P��yk�<�]�=-p~���l<�9�;��#>����k@�<(��<�>S`�W������P�^Y�V#�\���33� ʽ���<���:5`b�'�V<���<Do�=!��ȼXOȻp�R����e��.��=H�m�_��<W����)=���=��<��a<Җ����=��7�5W��[��13輱�o�,-p;��}����8�����W%���۩�^kǽ��'<i��`���Y˽Z��=L��:��=�-�=H��<�nr����3�<�[��?�������vκ���<]Y�=}�.�Z㽋���7���&W�����,�;�WP�[���F�=�T�=�=t˽�8=i��=,��=����5.����=�K�=��z�#���<�׽=�!>`�c o<�=��=>�������=PVN=%{C>:Y���3�<�f=��=@��<}xl�Q>�h�;�=��C�RP𼧃�<�x���6�޴��N[K=v��=) �;�T�=���B:
�W=��=���=R�N�0�8<��=A�*>4d���P%=�g/=�L�=Ύ�����G�p���p����\<��9=e�0>��	����=^=b'>&9�
6�<	��=�m�=HxϽ�tY�0M��V���7=�R�=X�7����<U���#+="*���i=�>&�<"�M=B�=�	I>z&>}�*> �S>��3�i�z:l���*%�Y���9G)���u���;?��aN�*b�<�I�=���=G�">�E>2��;慫=���=��`��2�<�c�=�5�<��=�u�;+��}-�=6�X���R������<!�w�
��]1<a�j���[�cxԼ-�!=z>�=��=�=I=Ҷ=�o	>�=n��~�N=�K=������;�!��p��s�$�p���g~�������po= ��4���;W4��=N>sR>rb>�8>��=|Y�=�^>�l>��:�Z����BŽ�U�=�5���N(��M�X4'>C-I�\���@��/��Dս�4��|l��nٽ�L"�p὚V1�����O���V�;�P%��X��/���Z3�b�r��f'�<�U=��>�����T��|��=�1>=j4X���=�$�=�NF>^�<�x���=.I�=�I#<Vv�o���:�u�Q�y�g��*�����=��;�R*�N[�=�[=���=bQ^�o:N���ļ����cQ>� >�$>d{>m�i>y�8=�/Խ�_���9C>`g\=�����0�Q>F���T;�׏�Vk=��
�_}|����U��=���T��f���>�iʽ�C�<B��UT�=J�=�j�=T�wp�>�p?[6�=e5v��D�>��=(S�!�t��fq���S�g�a �>r�¿!C���8�?
�>PO>g�?u�>s�Y?h�W?/NνO�I=ՠZ?��O?e�?�=�>�'��B���V����3��Yƾ�Nپ*���5q,>m,p��c¾�ّ��:�>s�}�Y(���x`�ƞL?c�$?*�"?ɑ4?Z�P?��Z=̌1?>ɚ>�~[��|>`��=��>SJþ�:?6y�?Be_?�ߎ��»$?� �g�I��ay���,̿mݨ���=�������g/:�6x������ӏ>0�O?���>�?���?j���xQ?ӟ����T>�.�>F�<Q�N�Nn�QsA�{�ŽB��y;�&7y�����u�lO�=��>��*=�9۽
̼�3&�V���7��	��%eK�T�-���W�J&:���z�Ь�?�?Ӳ�?É�?;�U�)ġ:����P��?��9�����Qվ��>�	��>�*	�71�>8t��A�[���+ɽ΍�?N�?)��>��1?�?b��XZ�3f�j.��G���b����>��>�]�Upe�N�
�b(?��>&B�?8�B?��9=����S"��VϾ��=�v񼴕I>�Ľ�3����q��!{�>X=i�L����D��3��G>���>�zc�}X= ��>��?{X-><�y��/?iC�?�#�=z�H��I�>�:���y��q
�1����[e���=�2۾n��>ۯ�=ŕr���L?O?�O��������C��=�x�����=M��>
�(?|y�>��n=�h{?Nݵ?��G?yq��e�����f̾�&ÿ�
f��x�~�L^��y9?�嘼P=?��n?��?�ʽu��?�=�?H�?��?��=��?��=c{?�����9?#~;eD=>�)���>.�#��I>�I���;?���{?��K�:��4�>1)��	�=f��?�c���)��%?Q�?ѯM�4�=\�^=ֿn?p�C�l�پ�N��%Nx?�ʪ>7r(����=!?��=I�����N>�P����!�G�g�%���l�9��>�/�>Nވ>�m�>���>��8?EA��]<?��?;�>�F��=*?n/ ?�0*?�����<�����-�ݾ�h˾�a@��E\��<�������Q�_� �AI=��������*�=𘯽3})�L��?���?ݾT>(�@>s�^=���>�d�>���?�A?|�>tp�0�U?l����q��J�J�X�`+�B,	�:>���wԾ��#>���:9�>��TV.?�<g?�����ߌ�e �F`[>8��>�Pѿ��v��t>@����0>�`v��
�2��>�����H���>���ȅz���c���ܽ���f���`~���=@"R?�GY?x�h?���?yΙ>pu8=��$�/�>`.�=��I�$z�>�.N>�u��DxX��c����@>����,����R=��%��nL�񥺾�X��\x����,�0��ѽLi�=���'8�$�>�Is�hA�<�C?�-I�ņ!�{�������� Cξ�#3�pq{�q\?yF�X��>{9�?�?�S2>�i�>r�>�(�>_����ȿ}I���;?�9����{��q$���G��7l?q�~?��?CLI?�T;�s�=oʼH�=���C���j�����z��%A���=��~l��9>�Jʼ��D�n�>؂�?�^?�	��l��`I>^�>���>N�a��H�>����mu�>W8���U��&+o�G�a�?f��^�w�A��=�{������p��)�H���b>���cAE?Y�>���=���Vz?�n�?ӄ��&���ӾN����=�1>h}�?h��?Ɏ�<?��o8?Q�?�?n?�o>_7���+���f������m�ɽ�L�>8�����v>z��?�u?�J�>�>�j?�;?��{?]�����+�(W��z������>ʎ�=`$L�w�>=��R>�6��2����>��=��6��6G���ƽܨ>9A�� �f=4�����>{
.>U�������}w�>A�7��4����ߩ>Y�����.��I�����>��c��D!=/gy>�x������־�髽�(��`����?�O��� ���2�
��>�E?�>�@?L˻>�^I?�8?�JM>R3*>��(>���?��M?;����
���1�>MN޽�?K��>�Ɋ�)7���i`��KL�))>4(>Y~�=B5�>�z?h���> =?s�R�	<>j7�?R�����>%��?M�?�Ή?	��>�]?1k�aЉ=L&�> �u��y�)�?5�?���v۾�JP���켼6#?Z�?���>@�0?�g����˾�}���a�Y4��[g?s�X?�x����
�����P4�:}h?M�s>��2?��-��n>'�(��0>
��?m~_��T��K�>�%~?�:Ҿ� 8�5�ᾥ�R?�_�?��L��
�?͵5���ھ�#�ള>��o��z����?�`�>�0��/:'>�?�Z�?���0c����{���,��=T�4=�-y���>��?�/�?�<c?��[�ʥ/>2��>ܶc?�%?~�������㐿�A��
�=o�>�t�=O�Y� 4?���=���=[�%��?�	/?M������}J�����E�����u���}X���7=��ֽk����R?�_'?^>��>�\�>]yk?��=�^�?y,�?��>��=r�����=���<��7?����ڛB?��>P��=�h��p�T>w�?��}?�2�����{�G�P������k�ۼ��¾e�X�\x�>�X�>����=X>�,?��q>�ם<nCw��������=���������	��k�R'?��G?�b?9�e?l�><�����f?Z�E> !M?&�^?
�>�ӑ?@��>b!�{M��\�&��׽����g6P��6��0�u�ʫ2�E;������䩾?N�?��?1�0?4ɦ? �f����>&�ʾ6��ԙ>KT����G޾<��?���>�Dw?��;<����U�=�	�>��l�P����e]���N�5w=�#2���?����`w��R:���a;?Y=���*��h���_�>m˽�Ӣ�C��zo�*(�	ҩ��+a�xܝ�!QN?�v�uT�f�z?>�W��>��?��=?��>�E�>���>ݯ$>�c4�D�x�*�T�'��)�D�1���㼢���!�ÿz,��>���"��9բ���>���>���=�W��F8���9?�me�3Z��M�ý_|c?��?�r��Kc�����~��8�=���>2�>���>[	5>R�	�*S�?�Z-?�C����?�U�?���?�l�"�����q=������~?���p� �~L��o��{��MI�|�>5�?i?�ƶ>A2�>�Č=�b���x>VȠ��U?k2r?*����Lc��m���-{�>��m>������E?|�>O@�?�<�?RW>�Ե�u��=e�>�am�W�+����?�@[>�/4>�[��8Y�?3�?)�&?���=K�y�7���v��f�?�X�(���%���>`܂�����u��?�r-?y=�>��?�Ҳ?F�?6�m?,v<?U�?:� ?�����TI��0�N'��7��6I�2�;��'%�F_����U὾g&E��R�?gR�?h�?��?�W�=���>B4�> /B�>M??\�?ם:�P?rrq>|���J�E��[?{�?E��d	ӾVK��$9n?Ί|��X��Ȭ?�����>y��xR8>`���G�z;Ǿg<��r���$m�[N��E�=�"߾1->K%"=�=�>e)�? X>���>sm�>ǐK?ԑ�?_����=����>;�?tn޾%�I�ߤ{�f�Ӿ����1�Ph��s�.>�.c?:��Q��=Uc��1xC�������G?fg?�Y"=d~�>�?a(>bB��+�=�h��~N?�^,?���>�7?QB̾�A�>�7��5�=����>i�����>{*�0����_/�3}?�鷾�yM���ͽQE?#�ڙq�.��<��
@���>a��=�<?qw?$���^ƽ�&��'<?��2>���4\��0J��W���_E�V%���v�l�0?C=���W���"?L�/�M��>xT�>�k?\��?�Z�?�ɳ?�a?��?o��L¾�˾x�����0�2�࿋2����� ����>'�H�]��C/���/$����\��&ڿ��A?_b9?T��]h�?���>ad��*5`��`?�6j�.�e?�rd>ڶ�?o�5=s��?^�@�鱿�q >����tT�ҳо��k�Jl6�҉}���z�?j鿥#"�����o�n����ً��V��W<=߸�;�=R�?�?��>��>�@/?��?�hD>2ݎ�ˁ�"f�>���=�����ܿA70>��D?V� �"�׿���>6H�=�*=�~��;��K?qk���㻿�#����?V��?OW�!+��P	�?���?�h�?�Y�?�^�>x��@�~��T�?����X&��#^?�[r?樺�}Lm�[��#{�?���~Q쿏�ҿKW�?Y�?Aa� �@>���>��~��nP���}ܽN��x��:�?#����r#���_LE�WO)?�?~�F4h�=쉽J\	?��?�!�>#ῗ�鿸Ł�=�Ӽ�d��A�t��>�˖?�W?�S�s5Z>d<�u"���Ã?����^�?�+m�	���P����~>�-�0?`JȽA>�K����m?b%c��&����M��ђ����>$*�?��1?��ڿ:�=s��M���B�1�?��>�"�?s�.>,.~��Ε�J9g>"�x?��5��>���?
�<�ʓ>oc>�7�?N�=?^�j�Ԝ ���>ȣ��k�ۑ��[������O�=�+����ս�(;?Ӹ;�@�w?�ч�f�Z?�)�� �?��=S�>�~>?SJc�o��>�Ƃ?UbT>o?��?�c�?����A?(GG>��n?��Ҿ�r׽nV��}>d�пF����?z"?;v�?St����.��p��`��>u�������ҿ&��?�*��V�4��6\�c��?�V�>�R�>(�??��>�C�>޴�>h�+<L��>�#8?ʳ���8%"���X����)�ֿ�xA��_���?�S��C ��sc��'?׷6?�?�?�1t��ט�z,@o��=�����!�6��E�O>m�����8&w��3?��������P?clR��s�=\_�>E�v��O�\�>@��>a��?���?v��!?���?��U�fb�>R=r����u?����r�U�?'r��*��!0�T�Ͼ?�1��g��T�?��p��-Ծ����Jl�~���?Pﾮ���>F��.�>M9k?�|)=�As?���?L�f=���?j�=UD<1$�����>#�G�Uu"��-�>|s�������=C�=#A,����i>�/�?�F�?1:�?��
@ʧ���@�>J�?�r/@\%���"?��<X��?�=��R��o���e1x��
=?#�_?%�=&a?u�)>�C>��@N�V���q^�}|?r�f�M,��#繾-憿kFW?^�	�gO>��6�".E�y�u'�>a~?�<=Pי�ο��9ԣ>/�>X7t?�k�_`>L�?��!�w8>���<D�>ʞ����?�3��7/�>4�?�R�β��
_�>�k�?�f�?�z?h��?.�f�`���/�<Jd�z铽O����Qʾ�����پ]���96߿�J]��{?3R�+W?KI4?D���U��>eb�>`�?���ŖJ��Ľy�>1��?.��>���ҿ�&=�{x2���>R�ͼ����@����t(��Ӣ��Ҩ���y=^�M?�D(��������?T ?�?1�B[R��|�q�@�@��d�=�z>G����>w� ���=�?|�o?(�"��T|?c2�>^B�?��� >	�a���Y����?��۽W�?f�l?!�m?.������C_w?0�?��E?5�B>D"M?�n�=��*�͍����8��y	?��L��5�7��>�;�?Ё�![п�ֽ
fs>���խ2�꣼��If=<�<���٤1�J�ӽ�P�>;�i>�?ի�?�Cx��]`�`h�V�>��5��H��b���ΰ?6F�>��!�h�\��'?��"�F<��-z��'�>7?H�࿵�j>�dr��x(>��(�/^?I$�>�>�O��_[�W��>X�׿�Q�}(�S�ݾX��?l
�>���m�=�W&����?=�Ϳ������Qۿ�Y5�cg���֣�U��y��<a��<ܵ�>l(�F�0?�6c?;�?u�?�(P? ��?���?h%�?v�f?�~?ʣ�;�ܾ��?�O%�"|���s���0r�>�,I>�<�>?�@Am6?��@�j�?�B=����A����=�V >Aة�����6�>����?�P��p�z���?�?=>�s�d>���?#�?[�?��>���?h=�D�=�LI�o�J����#?^Ǩ��j����m?�?�?��!?��C>��?��=-(�>TC�>�K�?:�o>	�?�j�?���>��{��'~��<<N>D^�?��i���?A&Խ)��_[p>SC]?L=�?����� ��~P��B�?����)�����5L߿Kﾽ������*��D?>Q%о[��=���]�X�?N�?�oU�]�?)�;���<�A�.�?��+>9\⾹���3Y?4�?���>)�<�E5�?��?~�l?�;:��?���?pX@�>q?!,���Fz�9橿��"�X��G���c;���?@���
�d��">�5@ �������=��?��%��u���������,?�8?���;s��>EVF?�[Q?z�;n��1F���>�d���2�?C��?f�þ`wX?Qw�=9:-��]���+?gH?�8�?��k�H���=�/�ƿYq���=H�⻂3���X��c
�?'ŉ?Q
;����Q;����?�X=����2L���?�.�?�T�?�.F?8�~���?;��� S����s���?
�*�) ?/��Ӡ�>��B@˦����>-2?`8�d�rJ߾�����^>0늿LM񿏁�?{��> �(�D;N?j'?o>?~>>>I��>E���-�=��	>7j�<xN��#>�T�����������%?H}.���=P�?U@늿�ޓ�мn?q^?3]? ћ�	e�>*3X?:�>S�?誯<�i+=%ӿ��+�Y����q��W�<��0H�W�I>0�>�F?���y?����!�>F��>�5v?F�F�ζ�?��?�vA>�򝿖y>|PҾ_*�>�H�>�L�?��ھ�p�������E�>����p�X?{W����?�5�|`�=�ߠ�|�>�g:�F�u�YrC� +v�m�ÿ�N�>�֝>>� ?Q����)=���<s�:�=�a��B��|�?A�`?mV���t>f�j� >P?%�о�x>��>�\�o�~��-#�$u�뚿4\����u?ky?竑?N�?2���!��=�uO?���?����i�2?;:$@��D?0��\9U?d�)��^�?��b�D0��+E>^��>aN��O&�s�/>|R�>�/E����=���>ؚ�>�
 ��n�>k��?�(��N��?կ?�q0�Pk�?a,<?�-M?UU=6p�>[�P�/�>A����'+��ea?���>�A�?���Uռ?��h?'�?X�@?�_=Y?M��?��?>dI?���>pb�3��(b;el�̵>�/<Zsx>�ZL��j� �:��b��N\?�.��a�k�?qݽ/DX?����'�����>���a���?���nÄ�po�ad���>�˗���{>*��8��>�C?Wp9>��m�?�g��?���>lrp����?�D�����X?�Ľ7t ��S�? ٵ��a�>w2}��J�?�H?�V�?�ꉾ����p-?�@2�?DѺ?e��>�xA?�p�?Ob?�(���*��O:�>S��;iÀ?�)?nu�u��É==�x?��2?��j�ъ�=Q�>Rٺ?j0�����B᳿�b�?N��>�"�7\Կ�h0?�9P?��T#2��N?J#�M� ��IY>�J�<RR��I��<���]���Q��(��7�˾yE>D]�Hm��_�=*uF�Jo>Q��>l�?(��>�g?J�?�B*?/7I?��>މҽK���A�=
�(=���#��m>2���N���:�>G��������3��?L#]���G�%Ҁ>���>�(?s��>�?Z�?���]>&?�럽�r>�m�>=�?Q��CK?��?����1��+?IU�<Nk��`�򾟘���>��=���\X���>���>3	���m�zl�2u-����D�ח�|�@>��>Â�>m>a�:>��>��Z���^q���.��mƽ�������=h��>�M�>��_�*z<=k&�>܂�=���;t���F��p^�#�����g����4�c>��M�޼lH>�o?Q� ?��>r�?���>¢廵]Q�S���tiW�{*i�jžg7�t#����WyľQ酿��D�rc��?��,F>,�?Q\��m�>�)?`��eP^�nƮ>���=�(�<J$���~
��x��tļXaM�3>Ai?��Ͼ�W�K�	?��U>�J���n�2�þ�纼A�<)��&5{>��2��.+�jR�>Qx&>Yپ;��V��#����/)?��J?�5��7}<�A�>�>���"A?#l�=�pȽRZ����|�$���q�O ����՗d>�q��eq`����Tb߾�<���>�=�E<�ay��	�>�z���n>��?��8��y�=G9�>86?�4�OV?��>���K��9־�k �{-�n��Dd�������l��)� >w�=n 4?�p���j"�a?�>`�?���Y'�>y�1?�k�/2�\�?��O>#?�S#?�?���>���i�<����>��M>���=7F�>�h#?Ԕ��B���N�"�O�>�9�?b�?��U>�o�=Q�����^�>�1>��X�Xp�g�?r|e��s��x�>�K?���>XE?0>?W�?�L����>农���6�O
�=΢����־��?�W�f���;ɽ��>���/Ǿ�h>��]?x̮�z��>�?E�}?ĭ�<��=�M?�h=�'�ņ�;5��>�µ��R����Ѿ�C��_��%s쾐� �p���w��D����{�]~0��@�=>���� ��d>#%�>4<>[uĽ���?OG>
�`>�"�>m��>�"�lɸ>�
缁)!��Ʉ�3��	���y>_�q�о�f~<���Ȕ �)o�>.��V��>�?��6?���<� ���L?���==���3䟽is�<*����=i���NR��5�>GsU�|����p�i>6便����r�=�%�>@����{Q=��>��%?_��C?�D�>�
?n_߾�k>��m��� ?�&��A��E��Ρ������'��ʾ�j��/�C>�D���S
���>d\D�ww"��T���>+���瘾��>���>��h=؂x=¶>>�1?Mޓ=�`];}���{	����aɎ�Y�]�wN5�<tF>����C>�\�>Ű�>�?]�>��>3 =�Ez�給�pz4���_�I᫾�O�� 쾛����n����=�'�>�P?��>��>w+?'��=��Ch����>��6��m%����������� � ���f>嗷>8+�>�ڑ>y_�>��M?�	�=�a�>�H?DOH?^m.?��=����\̎>��>:Q�=�y��aؾLa�ȉ�R�=,R�^�Ѿk.��s��Tvb��]>���w��^-�Q�p�2���b6>�}!���>YA�>�����ξ����_�=��A>:��?���2�>�+2>�}?~6N���?G�=Vv��7C�y�ƾ���&����9,���j�RƐ>�.?�s?�Q�>]�>,O`?�ㆼ�Z?���vZ��
.o�@♾���vT����>_�W�_.>��=.�<�φ������L¾���=l��e$\�?�<�
?hJ뽷z?>���>�[>��=���<n�b<WO&=��x�@����t���6>"о!k���>;C�>g�=��>
1?7�(>B1X��\���`�>�W�w���I���.?��O������(�>p�2?KH�> 7?ra�>W�>�]=��9>�>���?J ޻�N�>u#�=�I�>����P�>�W��ơ�*�$�y��` ̾I��iZ��5�>�>i
w�D潪�Y>g��>rD?���>�['>~6�>�o?�ӽܮ^?�%;>�\M=�'>O����Q��Ί�wY.�q��X;��$D��qο�?*���>�x�>#v?�e!?���>�!?
�X=x~0�4n�E
j�ˡa>ex�Q��W:���e��+�e��=~ۇ<2�>Q�>Ԁ>7�o9�<B��>0]�>���<��>򐴾�K��m�>�mj>޾���v+�	@?n�:�N���^�J>Eq?4��\�����;b��>�k�����>��:?�&?Ÿ��l>`|:?R��| ����]l�&0�U"'�J�>9o�>��?e��>??o�??/�|>`]?*^u>���񚥽?�=��<ω!�1ڽ���=�
�?o���wN�>g��>��5?����V�?OY�=�Z\;�w���̪�Q�;N���N#�R��>�^?�w�>kd�=pV�>�L�>+�P?�7?�(�>�)?c�p?�$�?Gv9?�~�?g}:?ܵ�>�p��o��ph��H ?F�"����>���>"�K?�߽G&���$?�]>|w��� ��=��3�#�Ͼ`=��R4�Y� ���'���e>~c�>�cN����=���>��t=�
��*k���c��`�L��+�
�Ҿ���>�Ak�5, �j �+4	>�%U>J�!?�/�>��B�3u�>Z_�>�4X�_X,?-�<URJ����>�[�<�����W��UW�nC����о�Q��T ��T"��5���� ;�?�E>��ս�[�>��;��u�=�.?E��R�x>�L�>H �?ޮ����a?74?*����*�/1�>s��=o���'��`�Uˢ�����d��5G�4i(>���>�Wo��)D���?�vv>@�Ӿ%~
?��>K�����."�p2F�O��=�w>��4��X���ʽ��6>��A�>�L
��;�>�h�����w?�>3>�HK?Pz�� &��>�N>{�=����|�5۾%�</�=5���!>�O�z^�<�`<>T�[ST�H����>��$�>�d�>��#?��Y�_�=G3?�=�^�$Q�%��:�-����b�
�� ��猙=j*��`�3>���>�X�>Tm=�n���?�Wp���&���L���l�@e��0�>�2��r�>( ���>K|�ɾ�>ih5??����?�Q�>�>�>i�i>_��>��C>��>7 !�/mr�>羏�Y���վO]���2;��$9�� ���s<⊞>���>ӻB>6V�>y�=��>n�
��|�=���?'޽�M�=z�>��B?��ؽ
+?��c<����
侃��=3J���}L�6`4��+;�ϯ�C�=ZѾ��LվV��>c�?b�=V�<��>��->�{=TX'>l�>�@!>~�����=7yQ�υ�rЖ�N�脴�T�,��_��~=�|��ߙE=��w>+?�n?�*�>�??��i>��T���y>�>��?�!=���������=�O/>p��>�d��{>�m?�����#"�{6>��J>��.?��� ?��O>T��>��O����>i>>����M��\a���ѯ�_�"���۾�{���м�>����M{��I5�>�E?�s���=�}>W#>�,n��W����p=M��MI<��4%�?վ�=�>�G>����#�ғd���>!����6*>����r}�=� ��/�C>�)?�=�?`�>�P�>a��>8�B?��=��H���?k�)?�/�>�H�=�=	>�.�>pm��;�8��K��<�>^cX=p.�<(p���l�>�Ϗ<��L��x��o]�=}�����rJ�{?z̤�d��У���m>�徽B��}x��]�\�m����9�+N�֐��Q�S��=�4��^�=����C;{�j=�B�>ts?cN_?D��>Ӏ�>;�?_赼b%����Mo=��>��о~�z�\�Ҿ�D�R�[�B����4H?�2��)j�=�7�=��4?�AN=���>��P>VՃ?��H?�:?}�,?�"? �>��u?+�>�\���5�=[*/��D?�4j��&�>���q�>��澒,�=@D����M���Q�����ь�s��@#*��i���1?�_�?d�ɾ��$>�Ģ>��[>�b����=K�>��kV?vx�>$�>I�>�Y���C�tp��>a �-%��q�7;9�����_>(�4>N%;����E>�z]�d��d�h��JM���c���Pδ=�Ә�7F�G޽\�j=�37>��?��D?L_3?���>i�l���@���"�$#?A�D�-�˾�]�!4ֽ ���3z�˄m�.\��p�Ra#��N%����:�>
��>g��<�X��SE?����w�^�z+r�����e�� �-����Ut>��/�����]��`�?Tgt������۞�>F-=σ!�A�d�¦)�ۋ,�":=yd>��D��<EG���w>z!>J>?�"����=G ��h��%'=���>�Ϻ �Y={��3e=?Ƚ)_�<�u���w޾㌜�ξރ9���m��gy�����x���$?��>��=��">�׸>)����Ľ��=�ܪ�i
�>q�U>�+;?��E?����ش>�vn>b1[���(���L�4�W�ni��&�)��*$�[�O�J =��4վvо�0�=�@���2��<(:>3�.?u@�?l�>�%>�I�=M`�>�.�_��=D># Y��sV�|2?_d@?jR?M�>ܴL>�'�>W*�A���R+&?��׾ny�� ��R �z���ˤ�A}U>����5���E�+��?��Y�����Ⱦ��A?�ɷ;>X��5�?��F<v�?J9? S?��
?���>g�?K�?�6��"���nJ^��A�>	�Y�E雽��f��?�� >ˮ=>6c�+��>lm>�;_=HN�?9Q�?#W!��]4?DO�>2U���"�MY�>���>�8�> �6�����&w������0���"�qUI�œ��~!L�<h����,>|^]?"g���G�������>̿>06��8�->[$o�]�?�MW?���>W��ԗ���>t�����np�>U3������>m�����WB��㾯�?�CY�>�[��p�>?�;x? e?��=��&=���5���C><�Z���>ب��rg�=�*���;�;�?�O>��9��C?�9�>z.4�ã��d�>��T�b���U�
����>�">�>���>�%?���=A�>�&?kn�?Tv۾X��Jr���=F۾%����y�Ew�>�����߫<$�Ͼ��[��k�>j|>�Υ=���>�> Eh=���>�ŕ>�Ǭ�V�ݽ�"M>r��>
vh>C�T>%a?e??𹎾�]پ^�>��.þ_�>�u�>�]�>���k�=�.�=���>ُ?r�b?�,?x-5?�
?Z��'̓�='��!""�{�R>�ؐ=��	>Fa���Z>���;���Qռd�>6s?K�>#$�>�>�0?��m,�y�>>h[����'�>fc&�i�=�>w��\�Wg�>��?�?��>(�-?�t>�T?�q�=,�> �>:�=��;�X��f�H>y>�T�K;�q��[�A�taþ�h��l����������Nݩ��<�;�閼M"i=RK��tӽ�>Oɩ�&�ξ+�<����>�"m����>I.,?H�1?�?���=9?Q>���<���=+p[>���>,?Bo���'��p&�}X��A�;���>3�?[�?�q"�b��a��AH����!?��� ��CL?�L���+2��;���Ձ�%�n>���>^��=��=�?z�	8I���"����>���;]D����-��4�?��=M3>ي��w�Q?`��>�|>�z=��>"���'�Ľ2?�Hq>N��o�l>ړ7�;�(?�V�>���>���>A���i��^7�wn%?D�>��?��	=:�A?S=��>Y�>`��?�uI?��[?�)?�{?��>��-?j?��T?���>*5�>�=�5�>���<�R�>f��>�����g�b,Ǿ������b��e�!i�?j�?�p�?��J>�Fc?�;>?(�G?Ԝ�>)��=��>H�??򲓽$D�>�x�=/�s���I����+5�"z׾7��X���趎����<(����Ry�:y)���1>��>,Y�>}?�G�>����$��!��G�ſ���i�=�th;!���M>d?VM�4���v��Muɾ��o������(�C��h�s��U?:��AF��$ľ�>n��ąI<ϒ�I��>��ľm�=�5�>U�2?�!�W�=�&2?^�?��J��}W>��>�c�=��5���"?YR>�#>dܾH7𽨊��3.�8�M�v��=�ɇ?P�=?].�>�>W�$��=<��=$s>>p�b>dI�2&�J
+�n�d�a.��g�=��5?��>���X|�H�!>��>>��
���>�����Óc�)K��? ���׾8��%�4?$�?��>��?��=?�T�?�g�?t+s?A.n?�S�?�MT?.G�=��?���>�X?[��>H% ���\>��h?..�?���� ?�
?7	����'�$c�>a��>i��>�5(��O�=���>�m��$7�績ާ�� �ݾ4Tþz��>��]�m
��5U#=�6>:�=�aB�@k��r}��ý7�<���,�޲?0ߙ?}@�?�0j���=?�1L?��M?���=�J��f� �SG?���A�=�⽼����z޾�L,�����x`�Mn����Q�ɜ+��MþH`��yB�2�C�z1 �Wvw>f�>���B�=E��=��g?��>S%����>��"�-��> �;9��>�Id��ս|bI�����mï�j�ܾZ�B|��2$>S�=j�꾆�վ�M>#c ?Y����v>�ż=ݹ�n供�$>|M��n�W���;���XS?�h�?�_��oZ>&\?�l?&�G��D >��?���=
����K�>�8>�
.�g$�=�^	�3���4���ol����%Lc���M�8��?x~�x.Ƽ}�`�:v���=/��H��>��A��� �V;?�}f?>Y�>��[��`u�<;��_�>Q�8�G�B�� �:a.�+���T��8�R�Qr=w^?\;k?��>[�=�`)>�����e��*;"?`��>-���7���ܾ��þ�Ϥ��׽�����-��u�
BL���?=U����VC?ؽ8=�R��%���~�<AF�=�n��"��} ���eI�!+j�hx�����nýW$���
c�>k��>�dR���>���>��>��=m�>�A=��?τ�?�r\>�m�Ē>$)<���<�\�h� ?4?f>���<9/ɾG9���
��ߞ�9��$����1+=�7!> ��f��>MqT?���>_�T>�'?�^;>A��^��O��p>�B��C5��Ⱦwxq�;�|�rǀ���D�Bd>�8>R�'>�����/��vl>1Y?�.+?��-?��>n�>��?�	{?Ak�>f:A>	_G?k�3��\��|.=F�6�*Ǿ@^о���>� ��Fn��>E>�?��">,C�=y%"���|3��H�<���-�T�=�Oc��Wξn�>vC��[ަ�ӑ(���Y�ֱ(�@��=Zf�;fue�^�>n�þ:%�>��>���=O�t>/�^>�x������"��%�,�~��v��>�i?P���9���5R?Y��?�Xɽ�<^ii?@{>��=u�8>S흽=�>|�7?��>)jP?CF�>���>�e�>mW8�3j$�>M���^���������<\����c�W�w>�;���@_�����4�=>����!�䆳��3�>�����l���u�>��½�U���Lɽ).>�A�:��>�=e��Т��:��}�������tK=]G�<m���O���Κ=�A?=@�����k�=�x�=��=�D�>%]�>z�o>��ɼ�o>-Ԗ=)(N=e]=>��_�B��PM���y¾�?>�2���7�7}A>�MY�c���ճ�#�O>��<�K�=�cc�Z�=C�>���>>��=�>�>/�Z�o=�b������2Ľd�=��=�1u��Ӎغf�Խ�(>�����J��oX�8�';��������|���k��B�r}[=���=�?
b??-�M�ӳ�;�w�;Z>6|��b\>��G���2=���>���>���=�3�>��=��<����%=��v=Qy��=5���=G��>��\��Ƨ�F�Wt��߀@���7��?2>���� =��*�g#��r�8����=c�����Լ�>�/�>�I�>���>�>ž�ʾ.��s�<�vG�FI�{s����ͼ�]����2�7����IýҺ���wɾ8��>����?���>�N:>.�>I�i>����lIT<ɋ�=�_C>� >}\�=Y�/=u}_��EL�0��=+S>ؔF��	���8>3	�=M	�^j��a� �� ��4u>F�=>-4=���=�%>���=1�=��'����оi��䲾m�����>��>ϐ�<͋V=�"[<K4�>B�C��=��1;��[=�w~=t׈��g.���^�¾&����ED>ׯT>��ՌV����<[���?���i=>�o=�{�=�Bڽ�m�]>Z�=��)�腚>[��=�Z�>�篽(�`=s~�=��>m0Ӽ�A�����Zg�W����z��M�������E���Ό=�3������)�o�>FP�>�f{��M���J>�F9>�{��T�>�1>���=#D�=��5>a^=׍���󯾚3>:k<�{>�#?����>|�����<P�E��F�冽ú�=���>P�+>m��=m�g����>�=6���&�#��>�.O>��>g�=�t�>�>濌>!�^>�4m>%�E��ｾoGɽ���>�2>܍���z�tJ>��p>y�r�G,��,�4>ÿ!>�P�=<3�vI�>h�=���> =�>���>�v�c�>�(8=�Q*=����Eý1B�B=������߾%�f�i举~�!��7�q��=R�>�@>��g=+ >pd����r���>>��2�r��=_͉=�|�>�q=�r���$�ތ7=Lb��$��` ������n�=������z�������澌K-���н��5�@�'>���NK�>^G�=��$>����b>9�$=��>��k�t�Ҽ�t���
�0s==O��'W�=T	�>�'�<�ע��h���hk>�|��t���\��[">v?�>���=t�T��>��>���=y�@>%��>�=>�iɽ�9��=�>2�@�S������<��_>^�����w(�ꊭ�B�>9=�=�+>G.�>�R�<T�ɽR�w�z��>�]�����L��Ǹ>��%>��?>��->ُ�>�<v�<2���Q,d=�ǔ��^�1"þMSb�,k��ہ=_r�=7���UR>���>N��>~w�>(ؿ<�D=,۽��=n�k[�ɥ1��HM��ٻ�46"<i�˽;���^8>���>��+>���>�S�=��>n�9>s�>}5Z��>�GpM����>�=�@�p\�B�=A?ߺ�>�v�>���>��G_��4�=�0}<�O�=�m�=��Q=�w��7��46���Խ �T�/l���Z���2&��,��~����e[H��m����=[3��{���
���(E�淏>��������3d����>6ԙ��v;+�;��\F�=���b��>�y�<�
�>��x>�Z�>g�q<�p�<�~�>���MY�� '�'���Y>�H.==��=���k�>��\>��^>� �=�>�����n=�}j>V��.�ƾ7̅��᩾�Nd>�d>[�=%�>�~4>�0��dU3��_<���>�L��d�t���=��><Ǜ<��=�WG>���=��d=-�����>�\�=�5�����?x�����>��|���-�G��<��>}*�=R=ۨ>n�=��A=�L��˼>=����Ƽt��o��>�C>O��=9�"[�>&L?Q��>���>��?�>@?�<��@>D�>$�?\jH>�^�>1�>y�>�7f�c�#=��>1�^��_��~����>[�"G>,�R>���=�Q>���=�&6>�D�=�k�>pr�-�>���>�G�>i������d��>  >5ad>��=�F��Z�;)Z=��<�P�<��R���%>��u>ڳ=��>���>"��>.��>M����#��SŽ���v���`/��|�k���𽔙�=��s��d���=��<��P�an��˻�=�(wp=�ۤ>�J��.u���-��:d>���]���󐾼v>�\	>�!<>���+>D��������7�ڼ�l�S;�>yk�=U6>�<S�tS->���=l�=�`޾����4��C��>�2�<1�>���<W]�>��>��>
O?�%�=��d�'7x=�{�>�xx����=��#"ἕ�ȽR�a>)
�=$o����>��>b�?�$"�X�>��=�p�>~H�����b���=)r\�wn�>A�>��?��>�a�>B�?ү�>&>?���>:�>��?�Ӽ>���>��#?tO?}>|_7�v
�F���a_�>��C��?�9>ˮ>�w��t��>C9��E�&>��K����<ϼ�d�|Sܾ��G��8G��M���j�~-�;���<�Zp�#7
�Y>���=}G�Hpx�wü⼨<i\��3��ג�>z��>�=��a��Ž�;���m�Ake>�<~���3���8=����O��yi��O��<&>1Ļ�8=�(�=~�_����=�@��ڵ�b!��r6�=��6�� ��?wJ>��=n�=�]j:\a��X����U��qm�=kxt>��T>V>�����gл�,>�}��;��/�k�ļ�IƾeR��Mk���9�N���-e�2%>��=��Z�He��s`>S�>̉t� 9\��D�>P���@[�wg��Dw�>��>������t�>��?����Z��>���=-�e>�Ǿ��>��j��=��>r�ܽNѩ��>�ټZ@*��a�����0�ʾ�<�+�g��*	�^ן�3,=~��=�y<pT����������2�>�7����>��0>J�u>�����S�>n?��>=�=(ʾ�0��m��4�Z���u���J�;~k�+��=ӡ��#��>��J>$�R>P�?��K�>�t�Ɛ-�Pd���й��|�4s��eh=U���<hؽ��>`�:�0@�=j�о$z�=��f�Az�=��绐[��ӗ>��J=�>�>�}R>��=�'�=�Z���>>J���E��z��59>�?>7� <%b���{g�>�\�=�_M>H��>*�Խn��>�\=D 뾴��>���>I�?~����0>��$>Z?�>(`�������Պ��H��;��r�p����IN�<�����0�߄>�?ce�=WK���	>�Β>�'�>�����9���Y}���=k�<_��_��h��By=�i;h�k��hB���%=@8�߬��ל�>t�>
�f>��>��>�&�>B��=N�=�<b���v����+�'>
i��^	�=�X��k>9�/�R�廩e�)��:'?=f�B�������=�`T>���>>L�s�����t<9��>�흾�ǜ�aվ����-����|ξ�5��#ý ր��os��{Y=�>�s����l=�4>T��=���<�4ؽDн�=/��n��CJ��q��e�I��Qc�G5*�\��=�� =�ᾀjq>� =(*>���£&>��G=u��a�>���>O�N>6�=Y�=�C�=�þr��m^%>HM�<w߷=�K�Kw">l�n�Օ�Ԯ+�p����)<�޽�V�Nk� ���W��qC���">���v垾�;����-=b�c��.�=�P,�,�=w�!�H�<z>��X��R��.���w�=�=vQ̽w�(��Y�=֗O>7w=��쓼���=��>=���=q����N�=�i	>�� >{N�W�=��j=�� >DH���ᖾ��Y������7������ʰǼ�
<�׃>$����|���K���>u�;wc���s���3>�7M>�)U>ގ�=R"�>N���=QL�����=5�c>��=��&o=��W>�E�="�������_6���=g�������Zk���"��o���B����⼴��<������9�Y�:�*5>R�u=�Gh���2�=��w=��x>l�=ۃ=+��>_J/��`��1�r�>=/[���0�R��f�����=F뽙/�=Fz�= �ռVި=⚡�v�=�K�9�2=��B��=��5=�) >:6ֽ��Y=Ț>��>�*�>d�>�#����N��ȶ^<�w�?ؽ030�@�����ν�5�0\��`3=�щ�E�x���]����>0B�>�PP>DA>p	z=�*�R����p�=Fz���W�#N<�}�=�(�=Q׵=�
=��>�|>�l�=6$<a��>�
<��>����K>`�`=���=�ͽ^0f> �<>]oR><��=w��=B���=��� ��e[�"Z�:�I>H�<��H��u�=
�h>�/>���2����u==�:$>(����/��$:�7!G�������x<�m=�r�<q�-�4m<I�h���=Ē:��'D��Ǽ<��/>��6��+�<���=�`=�U��W$>�R.>���=h1�
���̓�=yW>�G#��*�>�E���`������>k�ua���=j�3>��\=����(�=%�>`$>4���s�����=AA�=V�@�ؘ�>P)>���=
J>[�>�=�C#��D�<��>��p=0F�J����T>[�Q�p��{�'�C$>���=X->�&�>��<6���~b=ξ>!1S=�n<��%>a>�>���>�/�=I��=�E?)�4>�8	>6�<J��>{4�x������=�Z�>9�(�e�˽�7���T=>=��)�^�Y�?JQ>�Hm<>�>[�S>�8>�ӽ���=۞�<�'s>g8r���p=M=�=D�>��\����>�j���E:��ž�`ξ!����ѯ����J�� �Y�uz����Iċ��!=v7*�K���Ӫ�n K=�q�<�e=*�������}=�c�>V�н�V���s�w=}h�=�4���]��$���YTq��������u)>UB>O�6>@��P�=�Q�=?@�>�WA���&J�=�� >�~I���+�z�=��a<�:>L��.�>h�>��������<�潭�>�ṽ�As�lH�:�0>�P5=�Oۼ[��t�R>p�m ���8Q>��&>)ű<+\�=GH����4��t���2��R�8=�pi��뜾��{�����
>rt3=J��<L1>�2�;]t��b�8��Q�=k^��8�F�]��/>'4�=:��=��<��>����`�<�╽a��=�@
�dk)<���R�=p��:� >=�+;��EM==�>�lt>>��>{[��f�<��D�`b=��i��@��D�w��l�=Sm���=�e%�!9�=c��>C�>0E�>N��>�->��K�����Z�=n@�c;�O�H� ��=R�C=��G��"��=��>u>=j7�=Z>���=.L%=�r<[S��fa={>���=y�~����=�d�|<>㪧��֓�L�&�l��𺷾9Ӛ�T���O��ݮ�����o��c�9��E������O��=��4����+�1=���;��K<Ny˾q8���S����=�]���\��w=��G>�u�ۇ����Ͻ�K>��<|u����L�#���ʾ����<da���y�=;@�2=Ki�ooI=R� ���k�������H>Qxk�
��I�f�����4־�`>�[�"�`=>�=&->�r"�/�
�޽V>�B�<yئ<~�>#�\=%�K>���>��>Nx=*F�'�=��=�A��O� ʥ�8�O=ѿ#����z缝��>9z�=�o>��k>��%�WX"��@��[b>R�6�8���G�qA�>.W~=�[Ͻd�+���x>/ŕ>�[�>��y>���>��g<�ۼ7��=�c �E��=�r=�<E>�F�B� =�`�"��=!?üz묾����oc8ž�j�Xg�<�������D��=}2��$�:Y=�%�<B0?=V�2>�$=���i��(m<7>/=Q��b:=i�s�k�=B<}9�r���
�'=�O�=Y0�=ɼ�9J;"�>���>��>≶>�i��?��7��	-;�񢅽Ab�����<�}����	y�<gR��㒾X <�i��ׂ�(aľj�>�ѱ=��=��>�6��WNŽ���3�	>qp�=�o����<�JX>]_>><��<A#J�s�>��W����<N#�=��=Y�h�0|=Qu���g> *f�ʤ>����Z�=1r¾ܘ]��N8��e�j�>� >��>i��<J>�=�� >�y3>�=��z=���={�>p����$�Y����I�Ș�=�6>*��L�߾�]>�O�=���=�w�KO��q>+��=%ڃ���,�������ҽd~���k�=�>>Sn>�[	>��3>W�>�P�>!�=��>!u�>:m>�v">0�C>���>�t>C�C>�<�;�,>��=Y��>�w�\c>=ْ=c>>�.z��Ȼ$�T=zxC>=��<<<��ժ<D8>�ݗ�ePS���������BB��pֽ=q�=��`��>=}Y=�H�=bie��;˽2B��w}��Mp
�j�h�H�������p��=Y��d��<�c���E��G轗>�.��W5��Ij���Խb���X¥���&�p�콊��]���rӽ�ѽ�aZ�(	�<k�a�I�����:�'�e>-�>èP>�b>�Uݻ�<̶ݽ���+�=T�>�Q�<��6��>��,)I>6�>v㹾�M����q���s�V#��M��
������da�G>�=#�+2g��[S��>Q�>}�6�V�-�U6�=c	>��v�����ѼA�S�?Re;#㛾"��=f^=�0z>cB��@��= �;<A��>����Uk��[l����=}n�=�o[=�1><G>�˼���c��Q��=�׃���F<���co�=[Y��ϴ=��C<�Y뼨Ǻ��d����=�G=>�E����G9=?�E>Ⱥľj�⽤�2��K-><����8z�º����3�B<g��kɽ��=�;�>5*>��gi=���<.EW>��X�TZ�S
=T5=���� ���j ��hۈ�(!�=����<�R>��>�N>��%�}>o��=�P����=E١>HL�>�Wd>kh�>R�>Z�ѽ�������<6�>�v��
�R��o9>W�< C�<y7
�g�>���>��>�ߤ>�m�>B��=i	>��=����7�=�m>T�=�O��>��;o��=��>
���L[p�����n��'ƾ;Ʌ�7v��[����н�)�a��>)�>�G�=y��=&}�=���=R�	=�i��
�<?��=p��e������W˽�[�;_ki��n�/���˝=ۖ�<���=/��0;=5T�>t/�>*�>0�>�w�>�>��H=YN*>�(>2wM���o��[��U0J>��T��Xk�sݽ�>@_��X����&�����Y�=Eֽ\/�����2A>\�.�B{ľ(���X�=���=|������ǐ�mr��&���s?���ʽ7Έ����N���
R>��8>�d��=�=��>pƢ=y���L1_=#h'�v1��BF�Ɍ�t54���V�쾾/�	�zI�<��̼�\���C?=3>>���<D{��ڟ���་Ã�Uv�>)q�>>�>i��>~�M>��<4
�T\�=��>�U=�tC��&E��i�>T"=��۽^�a�����A�͗T��P���3q=���%I;�́�P
>9u��]��������>PE�=�<t����>Ii����!l?3��M�߾�`ҾES�>��?#����E>�Q?m���4�Q{��#�9?��?�O�ӧ�<K0�>����⊿�D?���>��?ڌ,=\վn�n=ٯ��ů������?���`]A?�Ŵ���_�&B:��)��l�����>ɭ�]��>B&.���*?�zT�c��>��U?��+���>��G�>?� ƾ��(@�о�??Lf�QTT=0���U~�͇�xfJ��?� &�q��<ʙp�̸�>G-Ⱦ��.xU����?��&?(r�RY���?����KB�#7�>�v�?Q�?&�r���Y?q�?h�&?��R>|�=�s=5$���|<��N?���%������]H?#�9?#?��F>����>S�=�6�Ρ쿀�E�!?�	?�6?�|?�K�?��лZs�?BK=?P�#?�q??�߼���*�>t!!��?�f�����=.?� ?~:�>KJ�>��?g��>�<l�߾��<�'�>0m���q?��뽪��J+���������=_��=\r?>u>!�|?;T��|6�=�>����ν�>����*�~��� ��Q�>+�=�ĉ?���Y���L΁>Ҿ5�㠄>^�>Q!{��j�?d-���K�>r���k��g��=�?CR4?_��rA2�����=Ea,��׶�8Y�?$��L��>#�
���?w�Ї��q��m�&?@��?Ӗ�?>��G1���� �k�����\?����\�z�?����ñ�/�>�'�>Da��%�=��z�����T:�����<w�<zO4�,�%�8�?_R���ֿ?�A>%�8��V;?�ֿ'�>چ�>˕�?�� ?`j>q����˞�8#���;�?����q?MrԾ0d�>�[4?�#?��=�!�>)�2?����N�&?�^	?f1�f ��=�qF�/����̿t�����Z��>�'%���?���O?Ĵ¿�J==��(���m��>[s]?4Q�>b>���f^I?P}�nu�>ǋ�># � �*�5?��ſ�*!���'?��ͼ���?���=W⿢���ʄ����*����!?Zx��z~><9���h�>��?������> "�>�!?Ăi���۾�5k�M���f��P�ſ8������=m1��K>�j��^K���)�;Ⱦ�ʌ>�ֻ>��(��������>�o쾲�{�f\>Iɾ�e�J6��~?�,���>R��>=7�>u��I���¾Г??��@�LL��5O=s�}�b�#≾�j�����w�X?� ���?��>�'[?�u���K�7����8�?� �>��3�).p��o?i߿9���������W?��/�&@�=�@���-��Cf>�H;<��>2��w�>�?�Fmc>=�T�=;}�>PѴ<�9���@����eȔ�t������\B�����k�>�] �&�'�n�¬�>��x�қJ>jqp>p �?�b�>c��?omW�R{��?���cn���b=�%U=Y=4�>$K���>�/�����.E�>K3!@3k����z�ǌ?��H�T9	��u�Nv+=�J��.�}Jw?�??��?��i?�8������?������>x?E>)߲�����DO���7�d  �	��>G@�<H�'�a>hޤ=�f%?�C�8=����#X�64.�@{�4��>q��>I�2?Vk�>���>��G?�?`� �!K�����>�/�?n��?���J��re�������K @? �O��?ʾo�E>Q%�KP�e�|����>�x=.������`�G;���?�􉿁J־��C���qq��}�P�6?9GC�Pv?��b>-��?�TX����;?�4�?�n_?2	K=ʧƾ�->�.x>���>���>�#��yV�1Z�����&_ÿ��&?EA��P�G��z�>�ϲ��ol>-�"?>6�?�/���eO>S ?���Y�����@���tj=U�}?��r>��?X��D?�Bv>2i>A+˾��>�����>$}⽃"�>hp9>�`�>�2f���?�>��)��Q�>��?"�>�	�>�R�>�pb�����p��>;?~?�~�>���?��>a�>Ub	>=��?^?�����}?���=[f#��W9�f���#���j�??tI?�ߣ?��>���D4?N�^u��~���q��?X�������2�P6n>��~�)��r	>�Z'�=�����qN���{�%�>�2?`��>�X��P�өQ�������?_�d?7�$����=�-n?e*��pt`�e��>���M#2�����H�d}??/�ϼ�"���n?r٦��䋿��v��;�<g5�>�K�>�D����>�A�=Ô��qӿ��%��	�B>��W�=���tG>�˾���utB�}��?���?U��?�s�?��Y�ff���@�خ�>��W?��1?
豿�E'?ԽK�VQ#�^��d2�?��>E��*qx?�wd?�b��]<��?b����4?5]?�w<�>���L��ݍ?�?�M�
��T�M58��:%>&8x?/�+Q�?�>~�~8Y?EM�>�C���Y�U?�>�G>D:;𝇿*�ѾT����G��|̾����Ǹ�;��E�E޾>Jz���?�$����� ���w����׍���h��G�;�'��7|9��ʎ��� ��Q�>���>��Ѿ�f�����h ��*��C�c��m�<E�<N�̾��+��=��B�V�g?�>�� W���`�M?�p�?!b,�oݾ�TM�l�!�0i0?�Z�����٨@?������*�u�>���>���>Z�6?Pkn?��??O5�>��x?��C?��.?��p>xw&?��=?�]�>��#����>���?�$�d)?���s��F���?��?�����O�?�@�=&���=�Z�c���!�>�w����>���^P��~h)?��~>	
���6�{o�>)�?�љ?�`?�l�?��K?]��>�:�>o}I�S�Q����?�J��mo���>!v?�ֈ?z?�%���w����L��Z�"�=T�? �ۿ��1?Y��<y#x=1�L�g|�>��q��B�?A�潵����䨿B��!W����F��{ƿ�F�>��?�������&�>f���ͦ��ӿ;�L?�`u?�W�>E�c�kZ�;��Hƽ�2���"�����h�?{�¾c��`I��ാ��Q�d= `'>&�0� ,I�!�?6 ��h\?;�п�Z߾'?���nF;���>xt!>O���۩C�lBo?��>G�	?Ϫ�!��>��~�� M�����L޿�� ?�b���'?�J���.=N��>@zt�͏�?"��X�O?a��$u����O�l>��)�
X�>�W�NNV?�X?�)_?j/7�z�i?i��_!>���b7�>-I�?^n�?�*���7l����r�C?#P?�)����?��*?������������'?�Gn?b��>s�������$E?�3����=�$V��Ww?A��=<DI?v�r���?��A��̕�,`��i�<����FCc��it�@2���i����>��`��� �{oٺ����Y��>��?��(>���>���+f��	ρ�	2y=N�bB����>�g�`?��G?�T��b���˿x��>��Ž����*�>'�> �=��M?���?���>��_>�h����;?V�>6<D��L�?cr-?!,(�5e[?�3=?b%ݾ�>ڃ�>z������=4"�r��?x1&��/?�>>������?/<�>ɳ1<.	'>�yɿQe+�w��9 >��?]Cj�+!���l�>�&??�>���>p����ȯ�j�7?>�Y�rR�>��=��C>.�Y�@�������Q'
?��r��1}�𦜾�=t1P?(̞��(Y>9�ɾ�k��$��>W>��>��>��?��N��A��&f?W&Ӿџ����T�>�?̡�?/La��>�����ܯ>���?z=�Q����{����?�e?β�?�wӾ�N>�l>iV@~a���~��8�=�� ?��>��=Á�<=œ?�6�XL�n#>e�>��l>ae?�?x"?dW�>6W*?���v�?.|g=�?�//=�9�>h >���>�Gu�M�>ԓ��3��A\?�X�>��?�eJ?pf[?F�=s�x?w���,(�5h{�%��>����4����SU�>��D��W��={7y>��~S��`�l>!��<��<<�>���>�
�?a g>S��>�O#>�Ƚ=�I�?��)�4ڥ>U�ȿk">p��>�F8��#��>���xO��뇽���Wy<؎t������>v��\���߾�d�b�ž�=�C�>\͇=^�L>0�� K�?I#�4?ྦྷ?f;?��?��Žf�+>�9�?>V�>ƾ�ǟ�_�X��_�>V%5��,�u���$��Z-��뺿["�>�P>q�?�r��|���V��;3�Sc�����眾]����|��N��_>N2�>�a�?I�3?R��;ʹl����=��p?�{A>�=��!:���a?x��>]����o��?�ۋ�#-���
�(��>��t�����$�f���+>�<�� ��v�>�y?4&�>���'?��3?uW�I�D�HϿ>�{>���3I:?��?6?��,�6��>u��>�MH?�e<�2�?Ȗվ%x+=��J�Xms?{�r?��νU��>�>D\$�.��=p�<�5��,?z"�N��Q�J>�!�>��B� Bk?uĚ�2�����>2f�>�
�Zv����	������ɾ�^����=���>
�>�c*>��=�A>	
��RZ�>�V>�+�>kU>?����ef�.1���w�>�禾W�D���(?��
>U(h�/2?n�?l�����+0�n��j���ɂ1?�??0���_�=�G��B�0?��U�?��Ծ�"�<����:�?�[<� &�?�I2>�*�>52"?�:>+������:�^�>9>Z�K?��H���>,a���� >j���M?��Ҿ#�S�ގ?�5]>Xܿ����R�]?���(�ĿcL��d�?�Fýp���˭=��?�x>fxS���>��>�i�~h�;	m����Ҿ�I�>��e���	��=~Ip?��?��p���t>5�3=�>D�=���?FK�>�V;��F�>�!�?��?Xa��:�־��!?]�9�[�9���Š>-
��=�_�4��D?�%�?���Y
4?����~��ߟ�� sV?vy�ig��܇>��U?����?�)>��y?B��>���?��=�oȿS��</O>��?:ÿ/�>j1�<`E>���Y#M�咡>��=����?�6��ڽ��\?C�u�D�ͽ /d�w��>��>�uW?�TX>��p>d<?���?��=v�>n0�?��$?y�;��@Q��0�?9P�<�\��`o���^A?��<>�z��鞎>�c1?���=�־S��9�(V?&���R�b�	�7�w�߿(s?������\�A���(�����냛��́���f���5> ��>��Y�=?�&?�]���>'�ʼ��M?k��y��w�=�:��o��C��E�L��\=<"�>FJ�<m'ž�s'�|��>�Ҿ�7��F?^�־�@�=e<-?�J"?Yҽ�8���n�>>k�������j��=��&��#�j>��d?�5�=�\7��5V>�V��U����?�u[�>�O>"�k?住��墽��W?S�F�䅿��=������Y���=~����9?x:(?{+�<����ҳ>��?�?�����㦾<��<�𻽀	?����=>��>�C���$
>D��>я�>%��Vu?yф�^���v��1f�>�;�>3�⾻J��o1�=Xѐ<HO�>>f���?�#��j}�>�E߾��6����wg�>��F?P�>�t�?�>�X���>�i?���>>8,>Wf���3���`��
�>��<b	l��-�=Y�>�F��>�
R��h�?Jb����~?[�<�݃���������c�>SG�?YC?���>5"?�Y�>c���BY9?�N!>��P]��w�?�|1>���<���",H?�+�>礓>~I>�T��j�=�p������ǀV�c|��a��K��>�v��+*L<�0���9L>7.Z����<��>M���^�G��9�>������>��Y���w��>�<Dn�=������>ګ�>&Ǿ����>;�A�QA�����?�)5��}־Rs�>u��>�'2��S?~�>!ľK[�!��=��:����4���������f����큾!�=rn�>�W�>V�=?+Mv�%�>[��>�>(�'=�>�s� ����킿��7��KS>g���1��<������>*�ľ�~�>B?4?(@?ly����B�JH>�J�Hx�=�?"|��m>l'����)?�KJ?�{���=�֤>��>b�6��{q>\r��t� >8�r�o��K�Y���ѽ,8����k�=���>���=�K�Ծ�0�>��}��֊�v�T>Q��=��	�x��;JE?k��?ǯ�f4 ��8��3? 5�T]C����==��>gk�>m�>��?�=�=̆8��\��Ԣ�>&���=��ۄ�<���{��?G����^�>ͬ���2���.95?���K̥�#�M�[�i?�Ӹ=E���!>p�?a������>6��x=?P�>��^��	v��5�>X�Y?�J=ֺ��sĮ>
N3?�oa?O$��H����>.~�>W9?�Z�?MQ?�b:��S��#g��W	=���?l�k>]=Ͼ����?�����Ͼy(>"�_?g���X�C��١���2>�Se> �>mԽ=����˷
?|Ƌ?o/�>����p�?�n?=�V>z�?�b?�/�>�2b=��>ߖ6?�t��?�>���҉>�,�>3�!?�-���e=�,��(��?�E�-���H
�4'��) ?�?_x�>����ʐ?1?�?+��>�����>�-�>�A$?)Q� f�<�*?��>��O>�O$�`}?�P>�w�>C٢��	@��kG?�+Խ��E���>�I>+
�f���V���4=�!������G(��;�5��CԽhu?�5<K�$�M���� ���0?#?&�=�&Y���2�M��9�	�$:��@���?A*��rϽ��G>o�@�������<<;_����?���w[?2m^??�+?�m�?��A���<?��>ϓ�>u�^����=pkq��>�?-�?�C�>O>m����>�'G�O#\>��>���>��1?v��> �2�@h�?"�>>;>�? 쁾䬼>�,{�ĳ;?��)?�.����>"��=&k���??&�羮.:�-��~��=[$=��?�Ґ>l� ?��B?�LF���)>Se3>�= ,	>}{I<�?�?&�?��˾t��=�/?M=�>�»>�ʎ��Q-?��־)J�> �>yr�>&20?3+?��;j�Q>���=� &�쐜=��ƽ�3��t�=���>�|?:̅��
��*�?�Ҁ?���=����⢽���?��'?�K>al>�"�?�P�>v�;�/�E?���?]��>)}����Z���?���.�x��P�|���9��.-��AŽ��*�,�=-�������>>����⃾�b���S?�=3�P?i�D�#��=�ș�?N�>�{>f��?�>l?VCx��)?���>|AQ>��>�>�q%�Q���_��Rb�z(����׾�}��-�=��?�Eu>��,?��8>�%�=��&����i�? �n~W?sdk�^f���->�X>�$<�}�>F	�>�\���W >�#��x���pPe�k1��E8��'z�=�(��l���=(?�*#�9��7C8?���=�(?ߛ�G �>�讼|�8�u»i�?�	���>�m��_Z?u�M��I�_>hE�@u]�ZV���}׾�C�?ם��Bx�,;.�y;)>�B��?Ož��*?��.�Dv>k6�DS[��������]�d>�����<�L;��q[��V��k�2=u��>r��?�5<��z�>�3?���ج
��I�7V��>hy�>$��b؞=���f�[����Η?p�/=�N?t⺾M%̿�@P�z���
?t���Z�?O�$?d�L���x�L?~q�������ʓ>>0=!��>Ŋ?�?�?��Z?ce����	?sV@勬><�1=�?Ɂ�>u"��>g�3?�m��Ծ�Nk��{���'���%��P?�Ww?�c���{?�p���_I?v�$>���4��ޭǽb�t?���=i�T���?�˿����W�?iX���[��C��
K�?]5A����?"Y�>&��?H�#��ˢ�.$?cۢ?��E�ȳX?�����_��ʁ��i?�%@�p%?�sW��2�>D�8?ȴ�2�K�H�ѿ���!��tZ�����>����!0���	?=�=���@cM��_"?���,��zK{��t�>?6f��r��8>�<�='�"��9�?��Z?L��>c�F=��?�F?�zȿ��l?��W<i	f�e�l����?��?��.? ��?9f��~����&*��"�>��G���?T��1�!�d�b�9��i��a���e�����M�߾F3?L%j=|�����>�P?�#2�!�M?-�m��q�>���>ʿ��i���=���=����K#?�i{�X��p�d=��#�{Ka?OG��U�=f1�=r^��x6���?�i�>i�����?tw	?��?O�>L���S�a>닅?�-ԼmAz?2^��i�?΋�>V�?Bj��<E� #W>$1ſ�K?�n�>��>�8��8y���I�N?�e�>��D?�c1������?�C �xD�������� ��r��>��?�R �E��>����A=���!r>1[�>���	��?��?��?�Y@?��4@#5^���>�̼�Ų�>1g1?�t*>�)�
P��!L�٭�>1�����=аY?�I�?�`5?�%	�^R���D?�����H�>Qu�>��T�>�>/?��-�&ew>�S'���c��0�e��>�C��h׺���N?�?�Q�><*��S��6O�?���?|�~���@?��?��?|CD>o~���6�=H�?}��>;���gC?s���t���J�>>��C�y�=�Q��je>@D�?�)���п>ݾ���#@?�O�������Q۽/�>��?�P*��W)=�c�>�?��U�t:3�=$��͖?���>�P<��*���'�<:�H�sJ�?��X>����:���?�?������G�]o���"�8,g�򬊿 ����Tb�É<��?��%����?%�>b/��#�'�Yr��Q>ɤ��e	���׈>�d�?a��h�N��U�{��=�_N�V��>�����~[?Fm??ݐ?�����|�??���?E�G?q+��O`"�c���p@���<��>=�?c���P/�����v�=�儿��{?����k�?����e��=���n?/���O�;-�K��?�q�?e;�?�ݱ?�"�>
����ܾ]g=�y��wS ���?D�?�X���/ھn�&�>�U=�m9���n?���W�	����յ�Ur
�����7?D񕺤a��%$Ϳ���?�Z�?�\A�D����\3>�J�>nش��ר�������;�0�ʾ�^�Q�F?(�ԽI���O�:>�s>
�?�������Z��q��Oi�*2ܿ́=���>v�?O���o/�#�?Yd�?p0?_���l����ľ14k��!��_j]?���>NTžf�g>�5&>�s�|DL?2�۾v�X�I+L>B~�?<w)��4�r���L�=i�?K�����"�lg?���3{?��a�$a??��/ǾцI?%����B�m���^l�� ��>,J�>^�?��S>7n��*��+M=��?(?�<�<Ͽ��?�Ȯ�]���#y>�1?�M�>�$�?`��>N�������@Jһ�k�J\J�?�f?�o?�P<j3@�����c��2w��iȿ��{?��W�sꇿow��?$@o��?D�m?��=�~M?�6��ʪu���
?�D>k[�<��={?�[�]�S�=k��?J+��c\��R��!o�>җ��ZA�C��>��s�!:>���=$�ƾT>�?��>��y�`����1��{�>S�$>����1
�JF�?��W�t1]�����"@?�&S��E>с�>�s�>����Y?AkM��5�#Ѿ-�?q������?�@.?�OW���j�˭��KZ`����3��>
1�>��*?\n��k�%�@D�>�}�>��=�>k�?�(�>���?�)>@N���}2��	��ʾ��-?Dl$�"nq?_1?�)@��M>�f/>�����@��8?�	��>˻�/׾(.9������H�>p�����?�8�?�Z?�W�3��g�����=��>߹y?��>�i��%g>��?��g?�3�?U��?ɣ�=,U�*�����>�%�>�>6r|?���"P?���?��?�E>0`?��[��K߾&a�=��j������F�?R�]��gd��'?!�?v"R���>�9��=�v>���0L�>����$�?F쓾$c?T�"?^9?�_5����?��?���>�*�(A?�;���=?�A���d?.��>�K��Ԧ?��?.žǧ?��?Ø���RX�ժ�{4x�"��>�S�?�+�?9������>�l��:VP���>���>?���
�-����?�_?��>{ؾ��?���>~��?�z������@H�?���������:N��R	�}�I>��� *�<~zD�ɉ?˴���C�?^�n=�ҽ����?S�?�G�)����Z��m�Z?�־���=?j�ǽ>.�?����>E?�פ��.�>bc�>a\>�I�ju>~��̌���>��G?5�\? ��>A`,?�:�?��D?Q�?���?Ĭ�?D�?�%�>RT�?R�?�dA�;�ʾ��g?�0>K��D�?�a�ތ>ȊJ�u��?�0����q���p?��k?�4r?�s��������>x���O+���	>#�g>�$��t�?	�n=Pz�>=[?��|a��B���d�?����g�4>Ί?>��,�2?l���~���nɿ�1����?A��4Q)?kN6?8�>b&��X��=ظ[>Ы����S���پ��>񴾑Ѿ�4�0ʾ(�ӿ����ޭ����k̾���>�����>nt@B� �����M?��>��>=ɿ���?")�=\�<4{�CT@���;p>bM�4�?� �����U��o�>[չ>�>?�����A���!?��a�¿C|�J=T8޾���?��v=I��>�0>0).���_?�W,?'!���+��ʶ�?W��>Ƭ ?�1A�S�]��ȿ����&�y�g�`~���e׿1�k@��?�%ο�[���[�?Q���(�?%j)����>cp�tp[��ys��}=���^ܾ�]�?=4���� �~-�?����V�=�??�fw?"�o���ӽ�D�>��>��n?��ྩN�ms>�Ž>�K���e������ݾ{�?��X����?U�x?Q���NϾ��p?�����H����I?^Q�>��g?�B����J��Π?��>��>��+�Ɨt>͕<�`�?���o-� �K�/���#*���?l������8�|�S$U�f�?&g@���?B{<?��>��=��@>�}6>�M�>u<��'?ż?�5:?<a8?��[�)��ˡ?��������Q߾r����P>�~����vܐ��N<�LW �(�^>�<?R
��� "?U�0��ʿm�M?آ��Th�GR4��$�<�k?82L�cLg����>#*��U�?�U?Io?Z�>i�\>`��>qV�=��1�pՋ��ݾI���k'�?o����>G�=�?�`��C���m̡?A�?;ͺ?�1[�zU�?��>	�?a �>l�>\�>��?�xR>��C���]?k���`n������Q�%�ɿ��?��6��� @[1��hg�?_��=��>�<d�l��>�� ?�����<�>ϨL?��=�j2?�>�>�=�ž��(�3��?�V�	ھ�j�?��?!��>�3�������T:?<�#��F��<���<��!��*a�>��>,A?��Ŀ���>٠>�
�?�;�=��>>O?}T��1�����>�>��>`s�=I�(���>��?��>t�K��Pi>b��Y�忽��>UÕ>}�>��b?��?��=�{U>aD?F�E>���>�?h��>?ȕ�Þ�gt������b�E�� ߿�h��݁�=��>�"˾��"> �>O�L��A���?�&�?_6b?��b?��+?���?�=���?��n�ϖ¾Zr>�<0?+�־E�ɾ�Ѓ>�R?)�>��œ���(�!E�������q�Y/�r/������$�]i�?��ؽ�H����;�b?���>��2@��̾�0&�y�7�\ޑ>��O=��g=����G��>�|>�ҾF	��=P�u��������B꾹�r=�]�%��=�>>L�3����������(�>�S>c��;!� �T��>4����p�����7��>�?�>�"?j��>��>>o��B�)X辢�����;9���������{9�;�;�����j�qiC��뀾��5�qN?��X��K?�o�>3���@�âl��O�>ri*?�K�>&�=�F�>b��>��>pW=��>.<��IG�;�A�>M�>�'F=�m>��M����>�#z>%=ν��t����>��龀G����_���>��+=XCS���0�4�߾�n��9�>�š�W������9�>6t?��>F��:O ���>�z��'�(H��w)�RRξx�-?�n�=�d�=4>5�-Δ����(��e���=Q���M�ET�>E@�5���P�?S�/=���<@����z>���6�����>�a�>a
�D���%U��[����F�����p����D������rC<���>��R��q.�_�E��{H?��?���T4��<��=������&��}?�b,??l>ɑg?m?����˂��8�=��J>��}>���;����t]>���>��b>dj����3�[��>�Hܽ�8?�
>�ڿ(�@��s*?q�d>� ʾX�>Klp?�W���R?5Q'?��/�g2�>�¾�8�> ��<��>lf�>�W;��X����>Tо�޾w. ?�M`�m�N�h��=��i��;#?}9T?s�[?Fa-������?B��?J3��4�^=�ZB?ǡ,?���� ��l*�+k��@,�����Wɘ������ ���?
��1���Ͼ��?�=�>�6�?"��iS�>g�>,�>��T>�۱?J�J��a�u�����۾!t�>~��>o�b?I���>�2��������A���j���k��t>��y>Yw ?:������
�>`? l�ʤ�=G�>g;�?Zȅ=�l�=H���׃�i_?9��;��>�A?_Ɨ>�
�u!V>�T3?��d<B׾�� >���>�+=q#9=���>�bi?
 �>�F�>u�!?\?. ԾO�L�	 ����>�T1;IO����	�������r����üB�->|�t��ݒ>-��>H[�#�i�ל>�Ӳ>��e�����z=��$>$Ή>�F�>T�8�ۉ"?���>
�s>�7f����:�'>P��> ^+�iL?���}����g��<(?~�>?c<?Mq?���?�w#�?�<�y����Ծ+"��0G=�ݼn��=X�JUY���/�?�1>���>U�>��C>~/���sv����=����l���Oʽ��0>	���i
A�<��EČ=��I>���>�t?Ǫ�><�p�YD?�ݴ?��V��>����R�&?�?�a?��1?�~���F>��@���D>K���������W����/�z�s� ��?>�5E�,��r�E>��a>i�w='�,>&XB=��1?:v���R���P�>KR�>�@�?���>�J>}݀?��ྥ�?��w?1<D?7v���ԾH���d��ؾ��=3Z潎[�?���>+&�����J�W��.���?HI�?	}F?�M�]z辽�I��Ј�hs���>���=I~u���:��=]j��
�3����Bᄾ\$�V�������[�>�v�_>��n>��?4�=���Pp¾�u]>l�P�\�ٽ(_�����%�j��=��@t�2�W>Mݾ��>_��>a��:��#���I"�C}�>���;�>��@�7w߾��m� �>��?{��>7�>kd,>k'?}C?�f�>��@h&c?�3�<�
���&?�[����H?9�?��?���־q�.��r�!�ľ�)�?��,>̱佬Qh=�4?H\>>$M�?!�,?��$��L�#!?��<c�
?�l�?z�J?� � �9>|P�>O��d)�(�>�C�=�Y3>&d�>c�6�|������?%t4?��??�8?.c-?�V�������D�ƽtA���)��Q����m����Ȅ�>�>̓�9��{��X>� ��&�Vz�IѼ>0X^�X�>z*}=�y�������?�\�>-O��%�'�]>���IT���=�Y>�*�p�>� �A�_?��^�y��$����gv>.�@�Q�t=�3?�U�>f�W�e�
��t����<�<�p>��?*��?��y?P���lm<���ˀ����>j��?5l?����]&�1��2������>E�?���>Ί��f ��{��>w-G=i�+���>�i(?���=-�K���`�:�T|v�H�l�Ƶ_?ɞK? <?�x?�ey?f�F?Q|#?r�>�3H?t>�?���?
�?���>� ?j$?@S&?���A*>���_�?�d��-,�������?&Y�� �>�m�st??
/��l���¾O����˾Ը#=((�J9��J��/$l>�Y�>�qt���=ܸ�>���>nN>V�=��X=��z�".��p!�?)C>�������*�<�<�>��2?Q���ʾ4�n��ys?���.*�>-
?J�,?�J���%�ҖP�4�㿈z�	#����E�о�[]��eT�\���_���|K=�Q�>�+>��T>�]>�������?Oc�������n�=�L?E���y�=9��>�B?����x�H�׼��=-d\<i\��ut=�B>v��	�����>۾�?�ݛ>'B��?90>�6�>Z����;L��>��=�C���.���b�<?f?��>�Ю������(>f8R=c��?w>���> 聽�D6?�B��+�>�o�E,�>N�T������j>rg�>�P�|�>4���+�>��>d3�>�P��F�>ht	=%���u���v>ɖk�ǚ>��<Bb�?cX��W�������>V����?�O�>'�h?9@��4^������K���ྈE>�c�>~��>�q��\ľw�����??<�<s�;>sŲ>Cn?c���(-y�&�q��}��H4_?���m�>e�>C,A>���=�\0?�����)�>�݌>\��>V����?i<?Q)/�"OJ?�X>@Q��+N����M>������Ⱦ��?����]�}���<�\�>k������>��T>��>��>J��?�t?~�9>=�Q�x
?�(��IN��<�?���?��@>��c�� �:p���Ծ�Dy��K�.I=�_��nӚ���&?�-�?�/m>z�H�����\I�=��>�:�=�{q�����[2P�VH��o�=�=y<@ҿ	��Lz�>�^2?�pE��3?� �������/?Q?$�"?�f?��Y?��*?���>�m����W=�D?}����z¿��;�^=�	��h�<�s���h��{������1�޾�����ב>���t��>�K�������ۊ�X'*>���-N?^��>��>�����;#/!>^ȡ��
̾�ڥ���}>��u�c��;l�=� ����=r���� o�������C[A��K��a��Sd�� ��C�>	4�=��!�q�)���>~���Y?��3�꒮�A4��ed���"�̿���T���X��j�F?��><p>[?�(�>��h�|W�� -?�<�<��ϻ2῾�ʾx�R����>���>�3��@�>:�$����������?��;(b�n���a�>���]����.�$�'?D�ؾ�氼63���9=�b=��o=�}->�Q=���hz�4ӊ�2Ž����H������(/>�u�=ބ�<e,G���>��>!;�>M�=3�>��(=�$=g�
���y=�_�=���=˅�=����C�˾\�*�	�W�hy�=��׽�}�I�>H�<��<�,=,��>4o=�=*�Q�нef�>VX�>A^�>VT�>z�>C�ѽ�Ϊ�)�Z��!@�=#5�=ɐ�=	���M@n>H�=��y>�󤾴��������F��+�ȾI���yۣ�Ôv��4Ӿ�Ќ=[�;��0>�ѩ����eod=�\\>&���q.>'�	���=?�>�>.
>�>��=�ڽ��n��˷=�J���`��G�`��=�L>��}�V�=E%�=4�>����lؼp�<m��<������pP>���=w.=�o���F�v��>1F�>�>��>üʾ]��m��+�=dO<�l�a���}��>>�b��ȵ���|�Zb������$����� ?j��>��w>��>qZ8=8�q=l/Ͻ�q�=m J<A T�I���3l�=K��==a
>V>�}P>u��=��X>���=�0B>
��=T���f�JX�=GR=�>A�R=�\	>SW>��U>Wy=�O�=R�����a�;����<���;!F��lCz���.>��|>Т�=	W�Xf��τ���<�5=��aʾ�`��XQ��+��͟�i�u��8W<�+���d4��.��I	=u�V��n����2xB�<2]���V+<7��=�Q���n�=~�<><�=`�c��0>hz2=��M>&֌�G$u���Ǿ�S����{��$����K��D�gľ�_��S(>*�H;�1�$�=T+m>�#>X����Ƚ�뒼�y�=�姾� �>Cv�>y$>2�>�{�>�� �|�=Ԡ��k�>�$�<k8��4�����>g�ʽ��=��(��7Z>�N>��>?�<�]�=hB�<��?a*7<��d��
'��h�>�<��=�W�=�(�>�b>��
>ղ*>.&�>9�T<^��~��<4t�>��@�,�@����Yz�>`;v;�ڌ<�1Y��9�>���d�B>�G=>��<>��p��>C;s>����_a4��~*>���=�!C��oL;$ou��vV;��o���;��#�b�ܾL<�@.�A��!񬾵��(8�N��=�Š�?��=ǆ<�T�޼��=K�>~�>>���6B���n=X(ս����&b���_7�=���Ϩ��g˾�샾Ѩ澧���i�L�>R�=��\>�4���=9�
=X9>�b���=T8�=G�z<������6�>�ʠd���>>���=(1>���>�x�GɽS�O�{->���r�贑�jz�>!!�>�-*>�t�<9��>܁E>5��>$5b>��`>�=O��:u=�D�5�</O�Zvȼ�m�"Ft>������Kғ�J��*��=��<�=�=���>�a�5T�/���J�=IꁾY�R!����=2 �=�Q'>a-~���>���=A㵽��Խ��0���<�寮�Z�<-�>�?�<y�ּ��s�*�-���>�ȣ>3Y�>�q�>��=�:&�ځ2�������p7��yNg�U��=��t�OS%�����!e�|��>��>��>_zr>	Q�=V,�=ub���,> |�D	�r�<d��>�(���۩�=� ��O��Jp�>�+�>Bu�>��>�>E>�s�=�$�>�h5>\�t=[�ܽ4s�<ҕU=I�0>�l�<_���>�R�h��l>���]�׾�*����G� .y��4�������½Osս�D�<������: �>��f|����C�=I�<�>,�	>�.>���Ž7�=���!�ɽEK¼Y�B;�ü�������������襾�C��8��<Y��<�Ğ�Z�K��qV=� ��i^���ʼ����w�=��=��Ӿ�����k�������>���=�H弭��=xO>�N����qᕼV
>�_�-&=ěk=i	�>��R>�l9>��S>��>��>)C�jX�<�1>(�U��e]�Gi�#o�<����G�=劺��>��}>��>�EA>q򈼗�`�4Ȏ���t>W�k�b���{[ =-D�>I�2=F*=�����=UNz>��>�2�>]x�>B$��u�<��:=@k�=ҝ�<7�1�_~=S�v��R���Qɼޚ�=�
U=�$�Ł��B'��J���W8���(�@��RW�����#��<���*T���&�=B)y�HT�%�׽��˽�|���I�=T�t���<�b�_�<���2�C���l=�l����2=�:9>�]�=�p�������>�-�>�X�>U�o>���w��+���	���A���-<��f+��V���*�������,}=�7��Q6�<ӡ�m����D����>]dq>j\T�륛>	�=�Ӹ�������>�k�����SF ��[�>��H>n�=W�<��>3.s���������(>(8^����=���<H��~�=��d=�D�=
 �����8r��EY���<�j>��g>�2)>�g!>��>�>'��=��M<S�)>���;d��=����?&Ľ2������<q�=OcQ�#;F;�ѕ:���Ũ�24>	E6=�\3>��N�
-y��n��R2��f��C �>���>�&9>��>�� ?��>Zʑ>]�;>�?}��>��>��3>���>];o>���>aa>U��Hp�<�>>fx�>�#:��@p>"e�=��>���[�h>�{3>��W>焛�pG�R���w �= ���Xl�D콣�y��xK�=�\�=�V���=�Y_>;�1�%@=���̩6�Q�V��[����"�#���+/�c姻�����B�=�W��R���;�Ui��]�
��6^��3�'6�������fFy=#4*��l+�~��(������Y^��+!��$�=H6�e`g��� ��d�>�+�=d�>��h�% ����="�������h�<���<)/�=�ʅ��.>�n=��>����y���[�� �Ƚ�~Ͼ}�þJן�bǹ�����t<X��;1�����*'>�y>�>K�{��d =n���#\�=�N��B���@G��'��im<����j��Y��ufC>p�о���:� B>ʆ�=V�����:�����	@�=�>�>�m7>�i!�8ս�fڽG���-^̽��A����>
1D=&q=|5�;U�3=�羋P ��wt�A0>�]���й=p�=�$>kH��������H<f�Ӽ�6ξ�W��ƾ{Ѹ�1ț�h��+�V��eI>�3��=%F<��=�B>j�X�q��=��3=]�μG��7�¾�n���5��24>o��=�}��@Ƚ�">w��=��*�ɃS=�FW>���=*C�=3q(>��>T��>�|�>#$�>�F=>�D��ԛ<�=��¼�D���o���<>h�<�	�����~n�=��>�E�> �>���>7ߋ=;"�>��{>��m�-{u=pi=W�>lѢ��J>��9�Hf>Kr������a���Bg���L���h1��y�	�z�X;$�1�ɽ�k�=$��=��Ƚ��=��>QP>m[�=��7�_�����$s>�^��
���X.���%�%�pNt���=�}�=u	��T?�-����>L�b>��2>D�>�K�>M�$>̑V>��=	�J>�N~�9���f����4K>��k��~\��(����u>�����Z���^��K2<ԕ�¯)=��	�hw�֌��% �lK�=*_�=����O��A+����¾��B��y;W��Vc��7]��jX��;��|��=$�>���4�=��e>_H*=.N>��k�����O��-<,�Ӿ�rh�}ZQ������d۾@��C�5�(�n湾\巽f�A=�r��k�U�i�}���{����>�>ˊ>$ގ>�q�>6�ƽ��M=�\⽹�>B�>$%���D�.��>A�Pa=Κ�<�.���Cƽ�9��Ho�=��g�󞹽�����1<����q��ɼN��>��U<jUe�Vּޠ�F�ؾ�Z>�1O�F�6>�"Y��Q�>h1�����Ӕ�=,��X�>Ϋ�=} ν�ݣ�	��=0W'?��?1��>��,?_g
?��	?Z�>���>O�'?�c%?��>.מּO����[3a��4�������������J�>[4_>���Y�>���>Q�������=�m[?8�1?���?��8?q*�?�2g?n�8�S>5?ɽ��>��I���!?+3��a�>(_X?��B?~
q�Q��=�[?ŔG>���]���i E�J�a�s+n�Y���P>�
?�ξ9����+���U?�C���}����>m��V�?�?���=51
>���>�=>�3������>��>����R�{�W�����V>�>ly�=�6��`5?ѝ>h?���ol�g�?}W��҉>R�>���;(�'��>��?�N�?*X�?�~�?(aW�F�^>�On�G���fp�c��=w0v�;)?���ޚZ=YwC�T$��	q����p�s���DҾ0�o?�4?\�Ⱦ8��;M)������/ >�վY��>���a=�~�.5���>Α`�,d�>7 Y>�X��>e?i����>�#`���"?�G'�xy�f��>���Z��>���>n���rՌ��L�>ԏ?ZY"���5�-�S�X�>���UѾ��H6˽��B?x�|�'"$?�?�>�i���K?����n���.����"�5�p��>h�>φ+=k�W=�[�zZ�>�M���>��>o`��-:?�O���3?9��C^�=��p�63�?i�Ⱦ]s���N>'W2?kVV>�q�]򎿑핿��h�m򼿩����9��>�Ɏ����>��+�gH2?[F��/���	��+��?g�&�ֻc�晣?�3�>L�0���?���>@3.?!��G?��=m�����f>�?�У>���差>wЮ?��(�?ޘu�z*��7r�>w�����?�g����>X�(���?I�:?�K?��n�>.��?NoU�E���£]>Ӿ�?{d�?�~�>#/?2�>].�by�>_�M�K��?_n�J?]8پ��?�0c>|���V�>���>�$�6�2?̵�?�7=\���;�?P��<�P?��7�?}�>G&?�x?��G����ǸǾ	�>�ϧ��[ҾԾr��5A����=�B�>8��J��[V.�̥���� �M��V)y>�ab� ff?�>�?�Tf��k�>�m��${�	�>sW�XAt;7�*?�����Y��$d��;����hn�=/��	6o�
;�>q�?�\>d;��m�'?e誽�Ԣ?����ӿ4?g�>>O�?�$�:��v�g1��I-?��%�
��>�13��F?E.��H���Ue�<��>�/�><�%��1_�wc�>��?q�߽Pą��_{>��B?��!?��>�B�>����Vؽ����A?y���R=���־8�`>w�ξ�Ю��{��R��*�= ˑ����>��>9\6�認���C�1��� w�4�#�!�u�8RY?���<�G��>*��=	[�`�'>��þ�T���t>p�����ʁ��#��Ѵ��Z0?�>�W>�i,>Lu�>�M$�������>qF�'	þ$��<�:����=�ٹ>ǌ ��$��y���>rG?�N_?�i?�2����Q>&�=�,H>U�?������o$?<Σ��=��-��*��`�?�f?
Q >�n}>���>��?�|�>���>�\N?<�:=���=P*>+��>Ƚ�>;��>����e���;�:�>��g>&=7��5������!#�>Ն >[M��}>���>���p�S�A����*W�c�i?�d8�a�1����=g�y?������?S?�b����o?֡�=4�T>�.�?�ʖ?�q���MB�3�#���@��N���>�mk>����2?��>O=��I��?T����{���?@VE?�r�{7&���O���M<�xB=kW�>񞝾�G���>��>E�N�p�+���O��=����.�<��P���8>I��=���>�ˍ�(>eЂ���:�;�=T�V>�:Ⱦ�b���=�=Ҝ>G���e�[�A�/���?���=��,�IҼ���<�g1�>`��W% ?���>�X����>N�e>�;���ھd5�>m��>�0$?9�-?^T?׼?�Ƿ<'��>�����?"�>yo=���;?=�9>ǤQ��7?tg?�b �GY��M�ʬ��w����0�!W?�r)�ӓ�>%&F�۠g?�jľ}��?k8?�'���`?�ί��-s>��j?��?�$��斾�H����>ka���,�G
���06�z�⾫��̮ľdþ�j�>%�P?*?�`u>��?Z4���C.��	���j^��E�>�-ɺ��b>+��dR�>V��Pɖ=��߾L������?w�O���(���;���?�H�<R��?[��r@t>y�A�\�P?ݟ�>ShV��x>�̐?F6ھ�9�����=/E�?O�C>|>�>��?��\������W?����?q����?�I�>��B?j����������b�>+8?\��qeC=�T?��">�
?'�>�Yν�5?|��?��4>�׆��RI�z)�Eܓ��1D?�
X�gc�>Ze\��+���m?�>X���B<?:W=�ר�>ӣ6��~1�G�r���w-��h0N>��>�7_>�?��*?Mu?�V*?
ݜ>	��?0a�>��h?��7?b��>��j?�P? �>���=(:�?IE>���)�%?k�a�"?��R�?�c�<t�<?��h��i�⤹� ��>��O���>�P�����1��"?�M������b����>C�>�{0>�� �s�̾ν�=�5���>�2�=�»����v�þ�
?�4��%�?v-�<�Y�G�/?�G5��;��b8�=�??=�7��g2=�Q�`)>ͧ��R'�G�����{�]��^(�tP`�Hď���D���?�?Ŷ?܇?T��?�.ξao�>�!;����=�@w>�S�>��#���4>��]?�k6?�Z-�6��P�;��|�k�x�{�=.��1�>Ü��ܡv?W���_e�?m+���5�2��>��}�3�Ͼ�R)>R�?��@?�}��T����&�_G?��V�:���F���>��g�윿h��׈��H��>���"N��Y��H�?�Y�=)h�7�?UN���/6>�zE�eY�>�Y~�q�ܾ�O>��o�@d�>G9��c'�􊄿�8�>���?A�s>M)e��d@��Z�?:g��?y�����+?q�)?|�?��=x�R� #)>�?��Z�O��=��G?�Nľ�Y����8?SD&�~��>^~g�[(O>�p?��@?yg ��qQ��h?�[���"���(�����>�	�>�� �" j?�׾�8>��+?V@?Y�O>�FS�X�<+�d��7�=�n>���y���q��/ᮾ"��Y?`��Zy�����>��ɺ���?����"-�>�p�?gU����?/V,�[`��>L�!>M���e�?���>��>���0J��$#�6�����I���	��~�>��b�쯻���j?l(=�=[^��>?���=+��>{u��%�=b!?��>DC1=�I��+!>���� Ѿ�#y�g�h� )v�$`�=r�#�-���^�^��a?lHt?e?.�?R�?@KN?p��>��?��2?�ʾ����_��>��>a� >�>����>z�?̡˾��h>���FK归]�>C�?]\���C>"O��𻸾���>:a>�q���'k>y������s&�=��'�7��"�!��
�=Ed�i�[�lҾ5@k?�]��m��>g�����>s�v=���>�ސ�$ѽ�?xG'>"��Ų����=A=>����xm?7q����9�-?.��>��Z�>J��CW�o��	�?�o�?HT2?ChB?��>6��>.�D�v�R�.Z?��\>%��>.�=o��=9Q0?BO=��e>� ���T?�4���,����=Yj?�	 �L#'��*��<?��V��/g=@x�� �??�Z2>W?>�OD� ���IG��n{��>���B��^�H�Ԃ�k{'��N?��H���S�=��y�7ƞ����S�;+���F>�.�>�<?%�V>�M�>���=�
y�1	e?ؘ�>!->�3�BC���̾�H������4�c���2��{d>}+��nf;Rw���(�>��K��~��>�<<�?� �>s��>��>��>���=�	��`�>�����\5?�V>��S>OM��$??{-(>���<Z>���i������;V���ξ���辽��a�q�����ԾSr^>�:8>I��^Vƾ�<d��.�=���-ˇ�p������?!�>���>�9>�=�ڨ>�>�"��!1+�>A=�
>V�ν1���}.>�^�>(V�=&쯽f]�>Z
�>[�8=-��ǫ��b>�v���=3��:L=�z�������|>��?��?Z�	?o/%?�9�y�߼.3p>c�^?����.p��^����e>:���:��=?<N<���9���d�y��<��P�^����>��>̳p>R�>p=�<T���Q>���8�}�j��
���M���:��U	��lԽ���=yM	�4�����=lQJ>Wy�\�B=" ��x\�?��=�j7�����GZ>��A3��oW�8	>�
����:������?�><�g>Kgc>�S�m]�>�>i 0��=ՠP>�s1>�z#�$�������l���Dܾ/Р=e�=�%�<8���Qȼ��`=�2��c9>M1$��?�|H=rb?��ὺآ=��>��v�9"-?�>�>�H�=�����sR?r>%>@@�=^	���s�K�����9ܾ����f��q���H����)>^�=���>������>�m�>�-w>ϰ�*N�>�.e>��=eOZ�W��>���>!}�>���=Qr�>9"���۽�A�;ݫ�=w|K<w������=�<�=F�^��&�BB��]r��>�A�=lH?	=�p�=�l^���?/I/�0������<s]�>��{�8>mep>֮?�	�>���>�y=� ?f[�����=t�j�Y`�>�I�b*�=���㫖>(Q��9��[>�F�>j���t�Q*�>(�>my9�&�>;��?@"�>3�R=#�?��?��>u�d�{�=�(���>\�ܾ/!�)J;Y��LK꾪,�<��=��(="�^57��:�>(�>����s@=۾Z?��>6{D>�>^]?��о�1�?;Ҿ<��K������G?�>�	b<�;���ھ�S@��������Sɾt����ʚ��qr>��yM����?���>�֘�̇)?q�M?�o�>c�]��34�N�̽�\ �~B=��>ȧ����>�R��=��h��EȞ=�Jp��>���S<\��>��=��>�U%>׌�>l�>�Ύ>��>��?w{(�%�>iy���U>������>�;kkK>>��Z���������E��=^�<Oa��Zb>R��O���O,	�&J>E|�������?��N%>%>>j3>o�����>��+>�Ǽ�<��rC�\n>��0���F�x�A�u��ꀯ��C/���=$��>>��>!�>Ij�>$�l>�&	����i�ܾ}f�=T&I�g�I=uL>��ؾ\ԫ��۽p7�>.��>� ?c7?WC3?�y5>�}�	��7{�=�3�Q�>���Q��X0>!4�D�ὖ���ݙ/>���>S�>��<��>#��Ƿ9�� x>��4?��@>�QA>�`�<�훽t&?��Z>���,�X����������ؾ�D����Ҿ�B���b���;ؾr��L��ũ��߾$�a0>H�=�m<����?��z>y�"�-^ξ��(�=�>*d?�Pe���?_
�=��=���>�I�>W�<9�T� � ����0ؾ�Z�����"��YSE>���>�Ic=wW7?F'�>��]=�"�>�U�>4��>:������󚾚9�����|I�>U-ǽs�[=9��=v�_>��޾Z����vV�q�,>
��T2����Q=���>> >p���8>�q�>��=�G=eO�o2�>yv�����I>�K��=���MUQ��z�=�Z�>Q�4>�h�<랃>�,�<�N�<�W�RI�>��/��#�	xa=�a�>�
��
=&�~=$�2?o�	?A�.?�;!?[3?�����="4�>ML#? �~�J�?@K��3�=jy�>35�>��c=dGY�f ���6����|"9���>��%>�e0>�5<K�u=��=^R�<�5?����e�?+K�>Aڼ �?�H?���>���	 �>{r4>|��=��s����>�����=���=�ɤ������(͘>�X?t\+?K?v?-5˾�;f��ﾖΌ��,ھP�I��2��C�Gᖾ�r�ܽ��Dx����L?���=̨Y��׾��;��>�4�=���>�H�	��@�;@��=�	)��x����*�'�{>CX�Qx|�p�=�W?�4@�CFV�~V۽��>���N�O���>x�>�]�v�>�N�>8z>�Ѿ7�6�	+'�'>b�|�2/6>�"�>�&�?�׫�E�?�#�=�
>�+�?�Do?@�m>g�C�:F=�]虾������3̧�oW=��;? �����?�{�=�`1>�?ܾ�:5?֕�<7��)�޾0�z�&o�������q��?��S?	w�>�8a?6~�>��>�^3?p*�>q�>	+?��?с?��?V�>uL�>Ҿ�>�3ž�����0�Yֲ>)%ľ�z��=�z?
!�>�^��4�?�K?��r>&� �r�>�𼶟��\#���U����K���`�j��<r6>�M���-��νd�>f���l��{����c��|�<��X���>HD=��޽O���r��U?�=�1=�`�>��t�{�T?�<H>�| �*
�>���> ��;g��\�>��>fZ��ǀ�p��>�{i�`�����r�����>�� ߺ;�Mv>	?���>�*�>��>�Y�a�Q����>��i�J?D�>4�z>�پ�;?2�=����s�ɾ� ��g��e��]�&ﺾK��������վ�����~Q�=�h�����>��r>�5!�t)�zy��x�}UF�ήu��2����	��Ua=T�=�n��f�Z<W�x���>�ɾٍ��̪I?f��=�'��{����>W�>���;���<�����G>�r�=���<o�&�X�޾�����H��C��Z>���Gh���꼧A>�v�|��EY����>�a�����c<�?P��>�����S?��w?�h�>?�4��7�ƶ/���#>�ھ�C���n��B�'>zʾa��2��?���>�����I?�A?%�~>�1�wԾ���#�>3�>����ƙ��Z��?*,���1>P����;�?�+�r%�5��>�j�0�C>U�<�7=)�Q=9�9Ξ]���<[Zj��սO
=Xh�>�����L��=[��>^��>6[?Ղ?��?�HH�:]�>�M�?�����?�#l>&<�1J�߭e?^U3>�@$�Q�߾�c��}\�l�H�@�羾����z���s{��:�=�;�<�J>rA<�(=>�]V<"�>�v�>ċM>\�����>c̑>� �=��@>ei�T��@��>�ՠ��,:�d =	ൾ�S	��z(�н>�l?:?}?q%3?�Ԕ>���> �>	H�<-:�>Qu3�� ��f+K�LI9>-Ã�Z��S	>��=�c��j��.���v">I��>,�k>h��v�?�N[=׀����VH�>_o��:��7�������:��}��ࣈ�����3g��Y�b�~:e�>��E�.�K�7��<`�> �=6�ѽb����O��<�;����Ͼ�?�4}m�͌��n���=7�=����y���
>I�?�;�:����z��>9?��R>��?��?�z�>sC>���>1P��˽�>r>A�?�)�=x�>��X>��>�'a>�Os��W�k��=�׿�O�k��ľ�*R>����,�F�߭��㾋<����K�qձ�hň?^$��)I��@l� À?7><��?S$۾Q�,���N���3�?�!��xb6�C�Wx̿P��ƿr�@4��Q��}������>?����bu?�����۾��}?�e�?�o?��̽�����>O�i>Â����9?}9��Y�>Įt>��<?�7��F¾�Y��8���1l��@��ƹ�>mD���?9?Si�>�`��[�(�C?�\?&�=F��q��?�~����?ꦾa�?�;>�(�>6R9���Q? ����V���}���	-�	5�0@ ?���?ެ@aKi�	��>�=h�p���Ͼk���<�?H�x7? ˚�oiO>�V�?�A?ow'���a��l����j>�P>#��=�$?�hJ?�T>A�p���S�z�?K�>|�ʻDS佔"�>�>E�	���j�?�%>3Cw>ƽ��v��-�>�T=Z1��V�L>2+%>�<�<]�?f�վ�ԾO��1
E?�o���'��ԛ�Mb�?Լg�90 �;}����?[͐?c*?$	�?�qd?޵P�3֑>���>-�;���>U9��p*�?����5r,?��?1�Y?��?u�?�F�?��{?Y��$����1����>L���>�s������^�ٽO���(p�>�Le������U��Qܾv�{?l�=y�?^���ѫ���>r$�?p!�?Π�=�@�w��<a�>-�����#?'XM��@^�aiھ�,��W�9?â�L��>1�?%�پ����E޾����cp?� B��3�>xſ���-�;E�mذ�o;�>N�b?�� ?v�?2~�>� ?<r ?3}�>y]����=�Lо��=S��=����ϻ�W~�?"��?V�>V�	@���>�H�����>��9�	[���B
�I����L��k���
���H�+"���>�:�?l܈?��D�>	�?�.��|a���L(�ltо����K��G;=>=vE��M��:��/�?d�e> ��>�Ӂ��8@�T�5�)�D�8�/��?�����&��ݓ��@��n?�q-?�a?�K�>"Q�T�A�i���j`F>��>X+�	�ſ��d?�E�>��>��>T�\�SV?���>i(�?:�s>Zt��[>��g؆?Ԥz����~߾��J?S�?F���ſf��ߦA?,�t��`��&c�x�Q���?�c�>�s>fb�?�3�E q?q�����A��ؾR���f�>���>8��B?�D�?ɾm�����=Q���S��HPs����>w N?�>/�?�(v����M�>ㅿjW�8y�?�h?B�`�Q���q��<k�L��Ф�|�۾c��??�о�R�=l'g>`S�?Z�X�z❾���=�r=d�&?�"x���Ͼ��3>�є>��_�!K�i�?��<���H�������?߭�?��?�2[?3�?H_�o���^o��B�����GM����h������>8Ɗ�����%��G�>�s#��6�?,a�>����:%��L�>���>�?$Iy���?���>I�/=E�6?�"?�F�>Z�#��ҕ�Q�?���>��ƾif>���O-�>� �>QY�?e�o?\�c?��s=:� ?Q�ȿH �1��>YB�?�ڿQѾ����H{�>���=�->�s? z��l�?�S?��F	?�{���憾�q��ҽq;'>��4?��˾(��>���=��Y?{3ؿ�yL�"��f	����>�)����?k��>��e?9[@�Ȑ?�-��z�ɽ�X$?��;?*�ÿ�$�X���"$?��ÿ������g?�L�>
>g8F�a��>��>}{�?Ÿ>����g��P[2?��?̂e?S�t>`��>�꙾R�l>;�ӿΪ���?��L<]CM>�[�>v^�>�	n�4�>۶?��N?z�'?��?��?���?q���y�(&����B�����}�o�򊚿��ȿ��O=���?��K>�\�>��w?�k�2d���:����j�
u�>��!?�?�>|Q۽�Z?��=>�=�=ڤ�����_F�>�Mj�ӕy�`3>���>9kV>�b�>^1?df�>�eD�h��>(Fh�T�>|��Z%ʿ�e��%93��K�����T�P���N?`�I? J�� ���>��
���?:�C?
ܼ����4�>��y?���*�?�?������?����mA?+��X�>V�>��,?�Y?�J���(Q?yXL�	]����\��9_=��@�wƾ�r���w	�(ء����x�{_�>�J@���>Tk)?�>m������S?��>�gd�?�퐿��c=٫�?��b?Ѿ����>�w�=��>En?3��>�6��iJ>7}S�����k�ǿP�>��?ζv>d�_?���>�G�=���?�%���2��W��?��H?>A���?#��>�m�? �ľ���>��d?G�g�T5�>�� ?@�ѿu	��W{���7?0�x�?ȕ��tz?D{�����u��=� ?��ֿ^��}���?�t�?|�?���*��z��?�?�V���?~&b��M?�����b��L�ut���y[����=�\?��}��/�'->[�о��?��4?��t?U�>���?^�v?��#?�d0�g�ҿƗ>�gF���}?a�l=X�>/w���Ŵ�,g>^��Q&�|�?^~�=�9?r �� w��WS�?-낾r�v>��Q��/�<��? �z�d=�n�>� @<�V??Mq>�sR<B�>/#�>9w=}�>�h�>V��>)�����<[���@>�d��p�?f+>|�)?pr�'G>s�?���>=�-��`���ӳ?�<����<���?E	�> ���q�V�?��z?Ź?��8=��?x�3?��>�/��t>Pp}>�p3�}ը?�8n?�����?�� ���?7�����u?�r?��Ѿ��>⾅�J���P��!��?�Ձ��*j>�e"�o@۽�Ȟ����?�\?pK!�7�̿�^q�1{��.�����꿕Q��U�Y??��=��J����?"5�֌A�<
u?��? �� �#>Z@�Ij�c�?q2�=��>��=a�<��I�0i��xԵ?)ݾ)x ?��?�go�X9�J]?�n�?g(�?5�y��1��@>g{8��'�>ٕԾ�鿬j�>�d$�S�
@����}t���K�=��^> .$��>����^?�r��J���
?9�@x�?��>�[?GWZ�h��%�鿈�Y?E0�?�>�o\���f�p�?�|>�¾P�ؿ0}���C�?7d���O���		���`�/m��6�E�
�"=;�<������x?X��?���ğ����#�>��>?����D��ՌI>�!4���>�E��0k>�W\�ق�?��u?�T@�U�Ӿ#,���I?̚�<�?>��������2���?�}ﾮ�8?_л�;o�>�{�=�ߝ�t�?�?�>k�>Ǎ/>:�T���Ǿ|�0�6�>���l�(�?r��}:����<��F�ho�>�f"@����,����> =/�w�>�x������>��%��Tw�?CX?F@I�[E*?<@��@�b9�?A�0��>��<>��s�Ї��в;�X����?�TW?@��?�5�>~p�>,3�?,��?�g�=x#���~?^�_�&��>��L�'�>@�o�@��>�a�h{}?���p?K�?§���?ꃂ�J�F��Mc?������>��d>u��=l.�y)���m��Y>��? GX>�q�?����>��s���]���P���C�����-�?z�?!�n>�A?�e�=rkP�e���jk���;ļ5?�]���H�?}u��QW�������e/�����Q�?���>B�Q��>N�z>ߢq?�C���׾�Џ?�����?1οr|���e��+��N`��]LF�O*f��K�6�>e��ʉ\?5QL���/����?���>;�s=�5?�����$�eU+?I���F.����d>�z�GH?z�>3�O?�JϾx�����+?@�3��1�>s]� �s�Z�����C?����~��Iſ�R�?=u�>��=�6ݾ�#>T�ܾ]1žA�����?�-?`ȿf ӿ���X���1��&>M��>��;��s�=�7��r�D>VF��df����?Ox�>��P�
^>î� �=3\�?8^>�j?�(Z��� ??Q	?����>WAC?�,�>�~/��7V�]����.)�%+���g�nE-�$�=�rY�p�>�*J�.�S>���>�vh�|����>���>���>~��>��?dŧ<Qϼ?+�6��*[��~�=!Ų���?J8��ƞ��HS?�$��(#b�>%����=f�����޽�*%�e���G�}�����c��u�?M� �Y�?��b��Q{?�?\?�<�@~8?��t?(���Y?>]��;��,�''>�T=�	Ŀ;����n��V�>���c��,R�=�k>?�eN��4�f8?`�������d]�JW����)?"��,�?��>����;�>�I�>1H�=�+�?{�J?=Ph?�0�?-e>����jX�>�ZZ?�'��5k?U ܾ�>���0�=�������>Ŭ
��E�<��Y����>�E;?G�D=1B�=���=2�,�׉�?��L?(%=
�B���5>�%�?"tս>�'�
�>�m={�?�~���>�����A���>'ک?\�?��?5���$����=܀�?y�n�>�S?�U��wy���[<�*?�/��w�-�"y�nQ>���?J�#?�d	@�=��@>���> �i>mM?h�x�����_<�3�Q�Ͼ�o� I�~?/gH=׀�=,(��3����1�J�;?�/,?W�����r���H=�v�?Nc>n~ >�ED? �5?�'�=#�`>��?��w?x�˽u�v�T������.N����=9���%�>q'�=�����;�z(>�(�>�%>g�v>Xm��P`�뽦*n�!��>5�l?����3�j>+�?O�7>c쪾�|�<(�P>��>E/���?j� ���$�s��B��>�rE>�����) �c�^���ӿ�dY�w�?�ꔿ�ȿ3�>	�?֑=��?�?#+?,��?0Zּݔ�?EW�?�;�?Vԙ��82��#?�9�@��>���>�>��@{��ysR�fo��,'=?�!�0��?x�>�?�>9�?�*��Ūg?}'�?P⍾Y^�i?��u?�%�?�����D/?}*_�`M?���-#��D}�TZ�=胙������C�mP½���S ��i?�*?�2��ŕ�?y�?��>�"��M�c���g?G����I?:.�?�Ŏ�#!��
�?
N���J��Is���`�Ͽ�I6�ڿ�acq��<`��.?	�>U~?�
?T��� 	ƾ5�?з�?�T >�5F���Y�4�g?&^S>t'"��.=nƎ�:>�Ѿo��n�$�q�>>�U��F*���A����2>y�K��>4�����>Ih'���`?fu�>rB$?��?��z?]ƒ?�{�?Ԥn��þ��H�~�>Z��sCw�r�g��??�>:��?�J�>rP?ƃ}��VR=ޏ �<�3�����=CI��B>��e���+��˙>P;�>c�	?����;� �>��?H��]��x�>�yw=GS��%wV���J����>�՗?�+s?{�S�L+��ž$��l��|�E?E�)?�����2?�-�<�A>>L���/��T?h��?'�>?�ܾ�:ǿ})(�>��>�&�>�x���)��_�J�6��!�Z��>��=�+>	��>  G�������c��#֐�j�>b!>Y_j=�I���P�M?�.�>wA'>*J�>80����	?�X2=��><�����>{��%�>v�_����%�)��^`�I��JȾ �W�24Q�Ѽ�>~X�=5�	!���{B>�q�?��L?4ƅ?o���Y��>*�?��@�m�?�S?i���[?�!�:��;>Cd��T��'�>�?E$��E澥� �E�J�$���ߕ?�=�z]?�{[>�,?XĿ? "?W�n=�!�j��>R�f?ほ<��=���=@���{ټTt���,�����g�=!|��G8��t���Y��VQ�8�3�9���R��>�I6���'p��d?�a޾�7����<m<?���=�۽t���c��>`X�+7>7���?(R�?�|?�L��ֲ�\QY?&o�>�kվ
��~ϩ>3G'?�3�����;�I�?����?o3?���>H"���>愆>T�>ɂ>J+7>��r<�U��C9�>�O?��?�aþ待��ǁ?]?+?k<�����I�� ƴ���%?�}==����?��½����3�?Xb ?j$�>��9?�6?Oi;>��h�A�;?��?��?�R5?�&��\���8{�>(T���E?��d�~BZn?+�����>���? �d?ֽ??���kR6�8�)���c<�Ɋ���x���X?�}�>TM�>F�>�>�^0?;��<��#?=T��;v#�eb��}ټ�� R�V��?�B�({�������(?��)�w#���-O��0�?���=I}n���B>�U�?囆>�������>�O�??��=�l�>^��>���?4�>/��<�PҾ5�=XǾ�=��1��|n�㾮?��x?O��=�P?����'���ҥ���	�=�?�>�^ʽz�ŽQk�>�w"���Y��r������ �����r�>Zv����=�x>�8?>�n���ؾ�d�?۵%?�b��v=zg�? ��v��?f>h7?�ʾ==��h?��?<�M>�I�>>3?]�A?�?�l�>kP��C~�>��>��8�����x��?��?ȀϾu~��sXF?�@�?G]��~�#������_�?Ŀ^�7���:�Ҏ1?6j�<H@+?bk>���M->>>�?9��>�p�>Vi>~�y?>y]?E��>Uվx��>Ֆ�>ʔ��V�?��f�>o��>c	�(�ž,ݕ����w�X?��p?�yg�ػ>&�ܾ����O��#��?=����8�����[���L>r�Q=7��*tv�q8>��Ⱦ��6��v���A>`�?���>yZ�>W����p�?.f��Zm=ܱP>X)B��Æ?Y3�>g3����>�@���x��p�?��>����[Ӿf��u�>��>-��Kd�g�T>�>W>e� ?�[���@��
?�?�y�}b���2���=H�s�b�9�5?��?���)HI����>F+�?��'�v>��m>��?H��A;�Íg���?��>�vR�FJ��
7=#�?�����?�=���2>�}ٽq;��?g�w��=��.��W@����Ĵ���>_�?�M�����>��
�I��>)���q�>�'T��8>Fy��L>�a�վ�#���L=*S_?�,���,�`�>���&=?�l	@���E�*>�j��To=͊-�״��b�.?=��_��<�p��<g��8���O���n�a�¾��=���<��{?]��L����X?ɤ�OҢ>�M@��F?Yµ>�ZԿk=)�b�����>��-?|;V���3��*����|>(�I?�l�>�>����?@Py9?� Ⱦ�d?Z"�=�}��g�Q����Q?TSH>��	��n��-@��h�4���R�+��#F=���h��=h!!>3���"?~�-?�t���*?#��=���>�5>��T?=XI>?Ɏ�b�\��6-?$��@7?�m\��bҾ[^? ��>�Bn���>5��>
�=�g?��>n�=��>����(�>�����:쟾��K�B�K�yPϾ��>_}%�J{���r>��?t�5=j}>!ݾ��L4J���@�nӿ]J??ݏ�>Dc��!?�(w>YM���_�?�:���^�=�N~?S�y��T���ҙ�����-�6�+����ν�����m�>�F�i�\>ޑ5?�ͽ�e����s�X�	>��?	�3���;��5���V���Xp��$��w5�L<Q?�j�>"(����%�A9?,���㎩����7�%��f�?�u�>w�K?c�j=:�=^!?��ӽ�Ơ�´}��Y��4��o��o��=��^����?�]�\U���m?�
)��O��l1�����?%�A?��Ͻi����� @�?O�W?H`���@���?c�>��I��~F��>Zd��L?�N>�,�>��>�0���R�>?7s���:������">����M�>�1?ِ%>���=A-�>�O��Y�M>J��=���Aq��s>b��>�T��E
�J����)��t+󾳔�� ����6�@q�>�s�>�ֽ��W=K>�O�>�!��{}y>�νmU>�B�>��>\�+<"m!?^�A�ܺB�)b�>D���"?�ꅅ>�����o˾�k���Tྒ�;�����C�<�K��+��j:�Cyþo����b����(�4>�h�����4����Y��a����C�hzh��{�=������B>ғ�>A���

>�?"�=]��� �14���>򾦽)��2�=:_���S��b��=�Ǉ>Yj=�?�>`��=l�̾�'>>O�>g�۾O�6=���=�e>����%(>:�P>��>H>"�Y��>�þ��y��j�>����<�>=~N�`��?1� �s�a�D�5?ǏB��M���P��J��ʂ�>��?��>��U��;>^[ �+�>�W�>uj��� ��.�uO���Ţ=}qh�6^>U�>�u=�挽�s^��ć>2g>?�D�=cm�>�#?\U��S%>\�>׃ھ-��=
��Im>lw"?��z?�J��m�'=��@>��I�N�>��<�/Ԩ�f�G�Rm@�B��s.�{w���p��$�U:�`�Py���QZ>ȃ)�]R+��ા�Ry>�"����B�־�p�"����j=�h�l�,>ђD��W�=q�=����h,�>�/4>�Dk���׾�
�>Z٫>`����V8>�!����پ��>�(A��z�B<}��� �����-�[��<��a=7?�t�=��=�?{�ξu:��2ip>h/�<t=�6D��"�&?ǭ> ?s,�>��>|U?�V=[�&��+�>30s>�G�>��U�c:?yl>��оV�-?��t>v�>ؤ>�<?��>��
?؜��BH�=��?�u>�|��-_+>o�>���>�P�>��>r(B>��1�Ȝ־Bs>����uѽ3g�>%�h>^��w]p?��_������؉?Qd0��^��^O>)VR<=U�=�2? <�>� ��Z��j#?�U�������0O?�P����ܽ��}�?!Kj�!�Y�B���i�x�A�p� <����\;�=Y��T���ھ>p�>�}��|��ݽ�>��:>����I�=Pж<�����!ý}�9<����tu��B~>Qɻ>���=o۲�#��=�6)�����$A��.��h��>�<����Gݙ> ��V��>�����>�B?����̾[�'���@��>��l>2n>g����>|{�>�(�>БQ>��>m>]~>���>��>�?�E���>	�=��"��\�\��>�N>�|����� ��Dd��0;�x5��3��%!�r�n���پP]������B}�;����i�T<js�?7�O>���翑>�%?$�:�h\�=G?��?�ю�2r��)�伢�z?)}�>�`�>�<��L�>�am>��k��1;?�	S>!��>��o����u�-�K�I�@M�=��]?:^?�t�>��>�Y���>���>��Ͼ�_^?��2��?�2�C� =^�z>�>��?�|�=�֩>�n�<?�=�R<>����	?O1=>�
�X���v*�P����G���'�*A�>y�?���>  ?խ����>��7>�|b����>q��=$�>�9�4��>���z!�|�O��xT<>�Z:>�9�>
%߾��}�*n���n�=M�Q>.���$D��ڮ�(8�o���4>��P>Q˺���C���>��>�?�T*>���>hq�>[��=M?
����+��V>���>N>����̒�P<��MѾ��ͽ�׸�F[�=D����z־�$�>�u�`Z�,+�Iu�>{J�=�DX=��<�6[�3Y��鍿�;8>/�d���\��>Ho�=�ھ��\�9[>V`>�Ծ�Д�f�=�!�>e�p>�(s>_��>V��ʬ
=y_M��ɵ>��=0X<��O?��?��E>�Q����@�]�3?�K�>cA�<I �?	�P����=��}���6>�V��X0�=fE=<�>D��V�">������Dq!�ep>�J��9�:a�˽l̫�(�	?>��-S�t�?0_U���7��! �h}s�>Q��	W���I5�W{�+.�̤��t���\��ߠ?����m,[��%���>�	��4� �
?W�;�� '��G	� ���/3>���=b�!>'�`�x���Mϰ��:�;zԞ�猉� P�¼�=y���,>.�>k�N>�5>c�U>k$�=�[��w`�h{�->��:���u��=��&���=.Nݾ� ��8�����^<�k�=���'��?�<0�����G?�x#?|���I�׾���>��?�G"�.?2�?��'>�����M��앾k�U?'����s��3�>{/�>�J����)�.?�u��G]�3ʞ���>ڗ�>=o=�$�(>Q���ғ2����>�/?1M?Ś轟t��=�\��sﾘݾ�Ҡ=��b>��>�>�'��`�x��񂾍�:�֡ ���?A��>W�Ͼ�kh>DZ�>0��um��Ej.?���OY=(��6�>kF$�ـ��"��V�>'�A?Z��>�">�؈>G��>��?�~�>߸"?%��>0�z>��>ة
?��>�]?�|�>N#�8�����C�K�r?K�3���(�{f��#D&?�=�����=-��>L��>��-���=��
>"�?���d�>+��>C��"=0�,?�U5?��=��N�>�>>�?Ok >t��R�>2��>�b�=5W
��k�CD�U�侂�;��P>��̾�)��kƽᓴ��=�>M�>�N�S��Ο���S�]��>9�����Nۃ����>�h�=w�6�+\�>�l�>��_>�C�<ǽ��K�>�/>���a&d?|�?.�=u�^�m����C��1>�:H?��辦�H����i��;?VH�<��>=4��>�)��D>"9�����hs=��v=����B�>�FM>Ʌc�୬����=�!K=�f�603��/�xkN��R�Ʊ��~�=o�K?�Տ�Ā+��?�u?�ֳ�r�-�-C?��>�؜��%S�x�.?rF=�>��8<�2���|�>N�N<)��>�3ؾ��1?7��=�i =�fa?U�>iH7?�>�j�=���
��=>�<�t=?ga�;YE���E�=\
�<.�7>=T�4��6��>�d���^��+�m=\�?��=��r�+���"�>�c|?�n�V9�=mU�?�z'�\K�b����?4N�>�*�7�>jS��JWо�vr>z^>-D��;�֊>�P�i�潎dB=�b?�yv>��c�>g�F?9�B?�\?%���6`>�hx=���>~���I�w?=Ge?p㗾v?���-��5��?��?��?�`>?9߶�J��>���>j�!�H S> �?6 l���>e�žߟ�>�oa>e8>�X�"����Ͼ"%>ֺ���[���Wt��\5�H��M�l�㏪�T��>e��>�X��UG�avɾ�=���󜖾��=7`j��Xm=t�=���>4��;�#	��O�?������s>.X&�/��>��>ͨ�>\�_?�(?1R=��>��>��>-�"����<%>/[2�-H@<�A�& I>�6�=�=о���>�ʌ>���J���`�G�RP �s�R<�ㆾu�t��I�=ANT�
�=�����*�e>!�ؾ,��Q���z(꾚�R�A�����b�Up(��~>������͌�P�e?����s�/�ʑ�>�y��>�ξ˰j��>��̾���JT��7��m!澛!���M��6꯾`_t><!�>^���~���=O(L? �׾3Ҿ6�?�?����>3*�>��+>Vρ>&�>LC?��?B�9��?B��>�b>�-���`=\�>)hs�Ǣ�>���>50�BL���CK�@�?�&��O1�#Ό�R"H?�s<M$������r?K��>���ټ����ς�Z�=���=[}u>�	�g�J�h�8�?=�[����3��JN>;�;#ê�x)�c8.=)�>���>I+j?�rz?�h>���>���>Š�=]
�>қ�>�#>����9�t;L���ʊ�w89��J����.��^ͽM�=���^� �=��뾲���w��U��>E��>v�Q>t�=u�>P�>��>Ta�>'�ڽ�F�=c�>�ZG��v��W�`>�ߧ>?a>@���x���2�ͫ�����tv��+k��=:v����1C�>s��>��p��tվs`>��>�?�ZǾ�g2�A�M>�kϼI'�>t}�=��=T_�>�l9>�o��O���"<J>٠�]�S���:�ܖ>�+Q<�/�=��><��=]�����'lV�~F=eg=7WF=FlW>]q%��µ��!��!>�~�> �?��>�d>�Tc�6�t�����?ؾf�\���X�%���W�>m ξ^��y���*Y��::߾�4 �5���	,ֽ��A>��I�U簼M{���/�������Ƚ.�=X��FV̾^�9���x�Ľ�=~�;>�ڼ��9�e����r���a>��R>n/�=,� �ž�d�
F�=��O=zp�>I��=i>R.��:׽o�>��>5���7��P�&_�>��>��V�ٙY�G�����<��e>u��>�ٽ;OȽ�G"���.��Ƒ�b!�xP;���b�k>��>0g�Qƾ���m>k�?M2�>F���<�B��k��`�>c�?}	�>2�U>�F>&P�=� >���<C�>�M�>=c>���3��I�L�$��v��⓽xy:=�b��Y���[p>�?>�,=[�(��y>+�v>;a�>0�%�6�5�g���
ܼ��̾T�?S��=�����=���>��)�-���t=�>xS����t��&�>w?� >9!��2��G�;A?=]v�=Z@=����"뙾��m����>Z������;pq��>��x� }?<�.>!%�>�O>�j��K#�u��>|�_� �=�y>���>p��η�� "��#�=fB����=�4�=|k>5v�|i`>��?�w>�����F>&�>�7>�&�?�{�vn>�%R={,�`e5�� �=P�'=Ü�Dʤ������s����
��K����9>��<!!�������=��?z�	�r�G�Q��=�谽�c?��>7Q?6{�>	=/>�,,;*���3�ļ09?1�=>�׾I�$�&u-�+����u���fZ��z7�1�ƾ�	?@�>L/�=�j�5;�u�<�,���af>qi�>���>1D^�l��w����^W��`�=��ڽGT��e =
|�����q���>�,��`q��A����>���=�Vƽ(��=rʤ>:��>���=��>�3?� ��OA���Wj<|uѽȵ[��ݯ��F�D����6���<�?Y�>ֽ��=�E�<*��nW�=d˽.���l�=<c��=[�޽�>V��k�G_�=�rm=�@=1t>D�>���>{������J����G>�h�=N��=�`�=~*�:���֭Y>e�>�"�>C��>.?���>�0�<�⾴P�6��鄏=vķ=�0ͽ���=�>���樾��)��mY>a��>���>�]v>���=J
>	^/������g�K���NE��{�=�Y�>{B�!�g��i>���>zD�>�Q�>kN�>�U�>�Ҽ��=�{
>�y>�5�:�US�wZ-��^<���=��k������r��1����*��H�̾o�о&/���T��>}�ʼ,�����[�l=ۏ�=�`�>	T������Ƴ���h��Q���(��x�>q�>]n'?��>��i�s��=�^6�m�=��>�<>�BS�.�� ��D0H�S5ɾ1���@@>\��>�c?鶇�ⶕ�Cbֺ����&ʽ���>�q> ���O��������E�p�"�>�A>2⡽�`��(D>f*ͼ�^���7��m>��,�* -�7�G��>��=\P>Yؚ>�t>('=w�3�����<�"��e��S��zc>��]�B%нCfA��1�>��=0�B>��]=�[�+Y���	��Og=��\�>���9{>���;�џ��"��st�=Ù�>c�>�->���=���=_�<I��>�,6?��)?'�]�oz�{�<��-dK=j&�>��>�k�G����#��9ó�� ��>~�(?F\���m�8,�=%h�>,�>�}k?S�
)p�q�`���D��;t����>�!B>��P��^r>�ؽ(���9���=��m�Z>���=� >U<�D	�>^?�?�+/?�u�>��>�D۾w���|B㾔�þL]�>��)�$9��v���;#w=o.��ˢ>�?����2�Ũ쾤���-��A��͜�=��:>��*>U3ǾH���f�����>�7�v�������s�>��zś���&>!�>��G�bR����}>�s�>���E>R%=��o=w��Æ�=�n�>�e>�������	��4�O��v�=��>Ն�>��>��[>�^>J�V>���<\P�<�+!>$�>�dν��ӓϽ7�=�S��j��>bwP?.�f?>Gk>-A=<ƥ]>��=���__�>)$?�z�>�$�*����F���~<�u�����>���>,��>g��>��E?�3R>���>�W�>��9?�^??V?��*?+��>P!�>
�>��>�� ���� ?i�>XP���j>��=���=��@�=��{>R$�>�8���_��!�=]�=V4����罊Cg�������ͽ5�9>1q�:z��ɽ�5&�y>�]׽�fg��"��T���ۣ�F�>��?�a5=����Rp�=9P�>c?GV^?��K�[��<�w���ʽA@𽹍�>t��=P ��H$�>$)־��]�b�=�����D�s[W��_�<m���R��.����?�-�>�m���y>�0?��>��>�&�7{�4=��+>�2>I��/~�=�Y�>��>^����)=���W��sž�HG�|,r���C�������<��>KU�=&�H�.@�)E�=��?>g&���i�=�|>O���O��Z�s뙼�t�> �=f$�L�����>?A?;Iž���<`X@����=�q��j�D��>�
?��p�ľ�2�=`�w>�>� �wlξ�E �G������=/J
>�\>���<�m�����q<>	b���tz<f�?�>'B�"*�=vM<�����+�JOo��_0>���>������>����)dp�ƣ"��d�����>c�>5i�g�&>��`=���i�u�L}<�ӳ>�J�>��¾�-�����=�H���4���\>��w>��d?�Y/�����Ӿ��>�j'<�R�>p��>��3>bu>Y2&>���>�K�>�D��u�h���(��}>ْ>=M+>yW<>m��>8����@�=R��=��>���>%�?�3�>�S�>	�?���> 28?����>�td>?d>۪���>~�?��>�O��:��2�Y������L���P�M�c>""@>. >f�=�-Y>nʞ=ØR=��<o�f>��?��?-�`�s9�n�����ƽYŗ=�n��HI ����\�3=�#�=/>���=*�w���|�q�ݽ}�G=��b>���>6�f>?e>���>QL=����ϯ=��">�^��HG���ˀ<g�>�k�)>�Rz.�
3�>�e�{�彤�ǽ1�?x
6>&�Z��%����=�B�=�i ����,�>H�c�
��;*���������(�Z= ��?!7��v�=dŐ��Z�*��KC>m&|=i��=<Sм�<�z�=8Ԣ<��<����<���3��(+�f���N�=���X5
�6���?��x=M�ݾ��l=�o��lV#�!�#��{�=�a<���>å�>TYw=���=���>�?/�8_��巼,�>J���������=�>a��</��2�=ĩ�>ɗ߽�� �ԟ����d>�_���XM�C�>qi�RD��+���i?d=>�Fc��VC���þ�j>���+���;>�{����;����
�>y6,�?
5�����b��>Í	�#��&��<��q��<XÎ?��>e��>��>�">�i�<�k}>�d?��h>�k� Z������Y�[d��9��>;w�I�
�y`>l{����E=�ǡ��%t>��Ǿ	^���	?(?S)4?G%>�DM>ƴ�>�e�>;RM;D@Ⱦ�_
�`��C=H��BS?o��=����˫>�I<�yU��p�M�>}�>O-T�Q� �]���3C>^���f�̽S�h?���#+��Ⱦ'j=�7\�Vn�=�I���]5>F����0?�E�>�;����ϑ>-r���`�XL�h�����>���y���&��
y=�*�B�<nm�>�s�//쾬����>�ܘ>.k�>����k�w�?�?r�#c���$%�:�>c��>�d�=�-L=em�U�>���}�n��^>z)A��G��:6�?�D���y%���P?u�s>=����\6�v�ͽf���.!�[\���L�=��>?�s>C�J��>;YX?�9�q6�>�>|G<��^e��>Z&�>�?���=��?"�>2�>�~=�_��Z�4��>����?  �����������>�(����XtH?*�Ծ)���<¥>U���<�?+�>N�K�L��4�=�k�>��>��K����,W�>��>
��@�<C��l��$�<UuT>Z�{��eƾZ���h�=����@�a>���=(����9t>�o=o�?�5�v���lu=m?>%�Y�"�	>��>�(��LA+?(�>D�����'�p�A��2�!I}�w흾B����J���N�G?5JN��\�>�@��a�b��6>��]���>bC]<UC�>"L��F7�� +>���c��=�Ї=$&�=;�Ӿ6/ ��$F�\G>qt;=ۆ�>x\��K V>����yj�In��m�>�B:?���>*{?��=��o>vn�U&s>���>?q��+�>�Y�>G�?�B����G}�>��8�j�a=%佾5>��?��>
��=��=�%����J>���>��=*�b?%����@���������T�=��f<�@?�b@�x�?lF+?��>�nٽ�S)���?N��>��P��(���?$q��Fb-�d����<����s��Ɲ<Ƿ��e�>�a��y���M�>>s�>���b�I�����oE>8�N>u)�>H��2��x��=�[�>RM?��{�Lf?�X?�ET�����?��V���!�r���s���	}=�L6?�R,?�!�����>�%1�в{?�m�~a>_j?�E�>乢�� >�ʒ�^ۍ>d�=s��\�>�?>;��>�-Q?�3>B�{�x���/l>�?:�J���?묾�X��K+=ҍ>���>��?�~_?��������UM���6�ϗ�>�O�>N��a�-�j쾅@��������>�a쾶��������~?ʤ�>��־PL��><z��#����=�Pa��眾�����a?f� =�:��AEy>@E���s(��:޽�97���>�d�>X)�>����&�����"��(KN���,?X�0=r!�>�/�>Q8���9O� �f���6��>�2O���>M=&�����Z�?�9	?T"?Ҙ	�>�>��%?Xk�>"y>��/�m��4���p��R<�9.�nMɺY��>ܯ��%��=�&>���h;��ei>��?O��>�:>?��fx��I6�>7q���}�>H��>ze?�$��&�ʈ!�W���k�#=�[J�����	>��>ֽ�>��>оwZ->������#>�>,>־$�=v��b_?+p:�u������;?q(5?ߑ]>��>\i�?s<�;�Y���`>�	b�D���=F�ͤ���Ҿ�F������+c���6d? �Ӽ��=��t?,4���ؽ�3����>�]>��}�|��iG����������?@��=FM(�8�)�4�>Q��7�Ͼ��ݾbe>4�����<#â��Z�>;�u�f٤��7=��D?��/><<7��<L��Y���h��8Ǿr�S<�9?�N��|��F,˾��;?��>���D?O�>D���:�����>)�4=4g׾牼����=��lՓ���$>@�?��?�>���>��>2D��nl[�/�?��M?��>�؎?_R�>
bU�ß���_>ά�=M�žT挾+��^h��Ļ�1	�>���>� �?�4:?��
�:�2���?�&?�\>�Zz?L���!�TT�At�>�㒾�%�I;{>}���W��bAk��'�>4��>��[�=3нG�>����C��=�V�>蛗>7?�?���>Zp�vIB�YT:�GP�������9�S
�>
��s���?��<�O=]��\���~�>e�V�g@����=op�Z ��@�?yFɽ�
��Z��H?��;�hv�>
��>���>����O�=��->L?��
<ʙ�Q�¾d"r?6@���X=p�^?4>ϙG=���z����?� �3ɍ�J8�>�XT�`tG��Cd���%?2?ⱷ>iBM?���O����V�L?���>���=\�Ҿ�G>�w5�&Ӿ�U�>&�?84�?����B`M�X�?���>լ���4?�~�>���<M�޾^-u��Hо�Un�z���5s��d�n?䚩?�v�?�>E�L?�:�?!h�?�%����>���?46?Ʒ_>p
M?�_�?$=>���=�8��wf>n�?�����w@���>��?(����K\�>�t�>*�6^����J=񥅾G'���>�>M<�R�	��='�c?#��=�yk�Z$=�d?���=:��ϋq>{Q<�i�K�վ��������=�z>��<?,�>�׏=�d1>�{���֘?EH��$y>�m�;4�a>D��>���=w��>����훿B2�MM��C�����&���>�DZ�Yf���U��;�> B�>��U��>�$�>�r����<a�ʽ�eA��0&?بs>)�
���=���>)>��S����X���>e=E
���ʺ��Lx����A>���=���<^;>�">ef���5>>�!�>~eR=_��>{�$��N?��4��iԾY�>�?��8L?�[ �k8>�; ?�q�?�����F>��,��,?�V�|���z�7?���'�z�1�Y��4G�}B�� �&>~?������O#ݾ�@��1>N�A>0W?7T�����> a��� �� �����r��w�G�>��y�$cT?�#��Xɾմ>~��>˥������A%�b���a{����^���ľ�]�?�Em�/3�;S�?��>W֢��Hɾ&��=ؽ�>���S�&>�Z��j����~>~�>��u=/���E[�:�>:K�>,Ӯ�v|N?�jڼg�s�6�?�A�>��?ԶF?��w>mQ=��G05��E����0O�>E6x>�'��8�>�������>�0�>�g�>u�N= ��>m�S�p�?d�?Ѳ>�s�=-�Q?�ƒ?��2�4?��>?��H�W���>pS�du(�?8��rm>S�R��>�3�>�O;R*?�9Ǽ�+�>�Ǽ��>q+2>y�;?d�>��j�b��>�_�=tk6�?���i)�}P*>���}ܒ?9,ҾV�"��W=3��:+}������RS?I�?&�T���=��>Ie��:��C�<P�>}������
���Ċ>r����e6�	�<��L>f�4�>�=A��w9>�)?��p>�O�=�">���=�?��Q:>,?W�F��d��<��P�� �����S> ��>/W?n�e>֔���T��?��4?�獽|��>�i�=�:V?-l���+�>X�l<�m�u��=�l�k%�/d���9�d����F>Ww�>O �>����｜9(�Y�1?�Q��,A����.?_����x:?�s>��E��=�>� Q�w���l ����>��s>D}�=�ɿ�w{>d�=�G���}�gE�>�
��q��,Ŀ��>l�}��|��-˿�#�>�c�O>�O]��V�?i��>膷�U��%㙼.��J������������>�Sm�3>?]�>ej>�����K���g�
�
?rN5?���>��м��ľ��?�\�?е&?]=?��q��Pg�7��?<?�t�=(��}J��v��,m^�BT��A�;=a���ϿfSݽ��Ϳ��> �1���>܊z��ѡ>�-�='�?�>��?-}2?{�?���t��?�p=�⌽���>?�[>�(�?UM>���<1�_�}��>c=<<�S�>��V�`@�>�"��T̚�0�=��,�5��߿�}>KJ�I��?$Xǿ�YZ�`G> ��?��	�z�׾_+�?G�����P?������Օ?,�Y=*�>��ȇ;T����T����Ӑh������U��CQ���E?p�>w��I�x��&��T0?MD����>+����� 6���	����>āi?ƥ�>�%d?sP?�;�Ta?�߯>��p?�]��ѥ����_���"?�+T��ھ�Ǥ��?W�R���r�fFm�*�?��e>D?�M>�g�<2�>(�׻�p�T�X=u��=�v?x�bf��w���9W��P3?.�!>R�?��r��E>�xj����>
�>�����??, ?i_�>jA{�aԖ=r����+?��?���?DL?|j��
��=N���W�-��G�><o��m*S?���=���>�?�?ˮǾ6��v�e�ޕ��:kn���������[�ɿ���;��_?���?;�;?�	������f>?S�L��b�p�?���>�X>?�y��T?հ�>X�Y�IH?�=�>��?2���??�-:>C*��F���ܾ�v.�X�Ŀ�#�8L��~���5����ؿ��><�?Tw7?���q�BIE?<�f?�}�g�?[!=c}?O���L�ڸ�!5�>��>�f���kz?��ǽLh��Y>��?-?�ڿ>��>�]��	�I���?·b�.���r�>r�?���5f�(K��g�@f*�����?ٹ���@:>�*>��;?6�?�%K?��?�v?:�P��'p�(ߔ�ޑ� �.?�^�>-��}��3"N?aY復��rGg�N�0>O�/�"/�<�D�>�9@��x�eԾ'4��V�y[��I�D��ֲ>�z��^���]��+�KW����y�`e���$���޼��#����N>V6e>N�|?�ݿY!�n��s��?*�	��]��]�?���H2?P�>���?�� ����>����V�MO�'n>>����@*�r����8>��BҊ���L�	�v�춋?���>�@1�����?Lb�d��D���l��7��>�辽eƿm���V';�0;���>Y����B˾�ă�=x��
�� ���.�>�����7���BϿt$?	�s�8>X�%>�=0?Ѳ�]�>��>&��?��f�����&��J�}��=�Jy�a��,;8�w�����+����U6���4���]��TO����>ص��!\����2?�:�c����d�������ʾ�z>�A��ӈ�匞�L�k>��>5�ؿ?�/?[��F;b�"%>�3@������w����?�h?I@n?t����Bj���>�\�с~;ĂĿ��0=,p�>Ȝ<��ྜྷ�:�^�q>mm�>���������y�.?Z?5?���>_�>\�<��`���?C��N����ž"�?(d��E!������/?Mz��1�d�f�=�)?2�?�l;?R<6>�/�>�n�!%>�<IG��v|>m�}?v芾���i��5�?��k��=�x���m�P�M��y�����7*�=V翼c2��,��M�?q����2?��>'?|	p=6B��n1ݽ��I���?*M�?�����>-�n��y�=*��>��	?��J=�F�l]k�q�ھ��J�5���r�ݺ�/<?��+?I��?�I�?䂃>�ߺ;�%��ԁ�?C��>���*ھ�Z�����=f�;��>��?�-���>�R���?�0���;b0��jf�"t���֩���X�KV����"�F��>��	?�zw��ן>�����>(�Ӿ��T�J�۾ԇ8;�����C�������>C̽A���1�>�?p^��T���
M>�d+?�L�>y�a�1�>p�-�2zs>g=i?H�9��ھ�J��yg�>�.ƾY�=�q >���?��?���=ˁ�=�z� ��>��M���T�5/�V��0�(���G��h
�S�ᾦe���j}?�¦?�\?�+��:A�<��??/�@4�X>�M@ %�(�?�n?�&�?s,1?���gdM����=�����2�{e>)���l�?I9��-�y�ja2��C�>�� ?-��>��Q?��?��>(�'���m�Z9���< ���?�ƻ>&�@>� ��{���ݐS?Rz�?��h>��)پ�3�?�İ��C�}'����>?)�?z>��=�ܿ���?G�����;?HWP��V�?��J�,�9>V�^?��?��\<���>I�#�݌>,���辅w$?U����=��b?�:?���=R���N�I�,�QO"������w�>X��?Z��?�>B>�?��?�+�>�N��|�>h.��o���S*��
����ri��!^D�PE�?Ԝ?8�н���?;�h�:?�?6���)5���g>�nl�]#]�k#�w@>��Y�Tz��.>�~�>d�	?����>�|�?��g?}�f?�?�2�?0\X?E�\?!30?���9؟>ATp�3쟾��$�+��b3�?P{��q5�>���>��྇1���s?G�>�v������YP��f�>�&4>�t��Cm;񶽾$_���8��]��<���᳽>l��>�]�>
��=P��=MM�>������.��29?`�?�H�?Ci>�-�=���>Z��?�q,�T�:���|?7�>���>�iw�>Fm��͝��q=>�!>0��ļ��<��ħ?h�v�v½�JN�Qd?|��=��>�խ>ߏ�?���?;�#?�y?�cf���?����3�Z�sy�=p��œ�?v��n]����=���=-qP>�-??`"�>�K��`��������>���>�U��(�=�i?�>�C{�T_E�[�?2�>��?b?�>Fy%>����=�=>��>��?��������P?�H�?RQt�
��>L�?�ŭ�����W>�L��+1��H�;����KRx�ٲ[=9� >�]i��LU?q�6?t����>��Ў��'$�	W%?�1?4x?[V����+��搾+��?Wa���^�g<�d7,�$.>�~n�?�/l>c���P�q�����uz��K=o�<s��>�lK��?n�>V�=#���*Q��:k��:�>�`~�.'�Πx>F���Ⱦ���>���>n��>��S�6? �K?5�<?�M�>�Z>1.)>�j=��k>�,��1Q?)Ώ�@�8?ܔ>cپ�}˽VN��nBL��*?Z�E?��
>�@�>�@o��ľ��we=��?���>ߩd?��[?�	+>��>�j@���?0[���?�%�xai?A����QL=�}i>�{�<���@@���9���r��X����C�dk;�1��=�o���W�:�v>�i�>f�
?�h�=�"?��?��>\bG>V6{?x�#>~��>D �C��9uɿV���-�?��=�	Z>@mʾѮ�?q!?dnK?�ٮ=� K?��}?k�|?.��?g	����F��m�>�b�>Mw9?5�>�_�>�7���۾ޓ���g�T6ֿcZ?���>�8�M�v>�º>��L>;u�?2��G��?�K*�������{�q86?��ؾ�$���Ŵ>H����y�W�K�G�˾^��*gF?�E���> J?=�?ۘk?]?�g�>٫?����Cp�o�]?T�o> �5��p-����\�t/Q?]N���@����M��?����� ���`9��K���X�1�[?Cߴ���>S�=�.9?�<*?Z�6>��?�
���T>�)�?�} �q�?�y鿚��r�>�A<��-ɽZ��?De$>�(��d4��Ɏ?��>O����= "?E�Q���ؾO��>N̼?I�>OW�W�@?p�>u�=��>q�=�9=�ʼ�� �f�F=��<�N�󒻽f*�=~͘<n���K��R�=΃(<���=	�,>$Ȅ=K�L��e�<���=e�6�W�=Ή}�}1m=����>����(��=���j�qő�����>YR�t���	n�j��=��S���<r��y�#>C��=m1,>��
>���>&�� ;��?Vf=�<��r/����>�	=����O(>��G=g�<=�Z����<����.D[�ӹ,�J�6���b�P�$����=���ų\=�}e=l¤=��m��1x��Ts=��W=sFD���z=ڴ�<[�=y6*>�	P>��=��S>pX=���j����==�
+�������@�I=�}�=t=�b<��q=I={���pf=L�»E��=�e��v��=F����ݳ=D�@��Ƚ�Rr=���=��>ek�>u��>���>~�D�7�=AB��]��K0�4���i�t�3=��:�j����&� �<����`z�=��l���]>�VW>��2>>@�>�ZJ��d.��{ۼ�5����@�u⽐����c�=R�c=z�Ͻ��ѿ�=t>>�@>ip�=��M=��y;�t�������Z=1M�=�ކ�lh�=��;��U=����UBq=�喾�P\����it��|_��=rUU��t��{	=�޼��H�4��<^�A<Ђ;f�<�r��^�~Q���?��C���{�=�5���~<MW�t;I�B��S��Ud�g,=w������=W(^�\��<ȵ<3�Խ���Ͽ�<��=��<�	)�đ=�����`�Y�L����l�]���������'������XX�(��)�m��O3=���:D���=N9>�I����e��<J�=j<��;�ȽUjG>�>g�\>5�=��{>B��Ϥ���j���>3@r����<v��-+r>;�=�>��37<�(�=>iM>w�=��>�WF=�͆=_�����>i%�!��<®�<���>�Oܽ�ia=MU>���>a
>�qP>�=��{>����= �<��I>�ح�#㛽���� >�b=�I=����fD>�ҽ��r>l3=>�c@>��2���#>s��=�G>�Q���׉>d
�>���=;4��KE�N�]����<FA(��5��-��T��o�X��X��a�I����6��Uq_=�$>��>��x��i�<�I$�C��=�t�=L>P���m?w���¼�R=�q̼�h���͘>�3��hu �{pB���k��rl��R��|u���j9��t�<��=�O	>.���W�=4��<��>UQ���M=��^<r��;7`D���5X�#}'�$3�=�c�=��>&P`>���=��@�����-�/>ē�v�@�͜��Q��=��O��=Y����=�r����S��C>A�>�m�R�C�d΄=��B=\����51��+�8�M�YT\��K��+���=c=�=�Q�='sd>kz�;�k�;�7�;�ߺ=�e��}��`p���=�V*>\�<����mG>M$H���K��w��AŬ=��/�R�A<P�ֽ�v=Z����P��R"=���<j%|>C�R>&*�>�/�>�tU��B�="	>ya�=X�E=M9�=�I�P�=+��6E{;##-=4��=�i�>lݼ>i'�>���>�po=�h����\=W�=��<�]7��#��R���H�k�K�F�)�n��;	-[>��;="B����=y4!<Z��<�>�;N� G���������%�:�H}�=\�����"�.��u�������G��1��괾I6��W�������C��v�z�lEǽ��)���ѽ��5��������U��Z|w���R��������J:�pr�;�"�wo4�@�
�[3a���mD��}u�={{<���� �辑9��"���ǰ�'�>�N�<Ƞ=(�|���G=a����Y>��<d�8>���=�R�=f3{=ܿZ�����U#�����Jt>*'n�s��=�L=��'>�
W�a�ɽ*�+�cW�=B��k�rM�<���>�牻�=r���=�]�>��ӽ�9�=��=J��=٫��c2��`��<��P�L�����F> ؈�D+��
�Q=�����DOŽ�DW=q��C���v[�`=@O�vh�=v=+P�<{�o>ق>�V<>���>87=P�d���VZ�͚F<1� ��=�n⽲��=(j�=�M��a۽��Fc��	����೾{4?=�ݶ<���8�]�y�=��<���=T��]�=C�<�%p=5���K=�{<��=���I�o��P:;̽�ƽ�� EV<�����-ļ�/L��+�V�<:.�=� p>�[�>�"}>���={����w���Ib� ��l��J@�h@7��KY��� � ,�<�ɽ�˪���6�#V��ԽDdi��=n)�=���}�v>�U|��X�đ���K>��؛)<�w~��H >�kb��<�=��y=���=�L��Զ)=�X������%���<�_�>�̐�I�'>a�<]�[=�[��B1�}��� ���#=��=��J>��=�'>�]�<_�P>�>q�>Ā>13�=��>�������� �Y�;g�����=��=i�m�E��^=��q<j���^t>vA�?R�=g)%�{6����[�k��QhG���>���=��>��`>��>mm�>馚>C�o>c��>[�>�0>��_>�M>X��>Z'>�r�=#�S�L<<H ��>��b�hZ�=��Ǽq�!>6+��Ǫ=+DS>���=AO���� d �3T=j"%��h�>�z� ���*�~�=�t<����-����=K7�=X:�<`|޽s;޼�ɼO��J�����=w'9���d��b�=Q�=�J�=,��=6n=����e�=c8�=�r�=��=
,=a��r#�=#�<{����;�@�=��R=��ǽe�����x���w0������u>p%�=I =���<E���g�<�(!=Pס��o<�_)>c�=Ԯ��H�r>m�=*
=oH�Ѻ���J��ʒ�b���k���k^������Ԍ���X<�@G>�r=��]�Ef<#��=2>�Dս�<�A�=�=�M+<�觾��:�Q��X�=���@=��=�5>�(��_��=�F=�V>G���ϼGs=y�u=��>Aʕ=�>+�>�4� ���
�=�<T;���ܠ<����6��=��:="����gٽd*=;䧾�H���=zc>|
���}=QvI=Ƀ$>��,���=���=H�>_�Y��8��mR��B���6����P���b=��[��=��t2���=�0��x=�=�,<�@�nmľ�6i�y���D��C/�:4p�>=(D�<6��ma;>aB�z��<�x��L�p=C<�<Ga>ߙ�=��>�>w�=O�==�m�=�M�=/5=j� <��|;[�N>�ڰ���=ms7=q�,>b�`>�[>���>��>�k�=:��=y22=Z�
�,�����=��<����]�>;���vͤ<�6���˽D�j�T����[�ؿ����6�;�����ν]��c��=/m�={�>6�<���==�&>ѵM>TUD�h�;��x>?K�=b��=�=Cb�<z
	= ��='=A>�x��7>�]=d�:o`�<�,>�>�%�>��>���>q��={��=��=�Ѻ(ř=��9|t�ڍ����=���Ja;wy���#>��=�`����$�z}�"���t
`��A���NN�����d����ܾoع<� �������S�G�4�t�%i5�����M��ZȽŃս�����-����<=�~>��=5�f=6�N>�}X>k� >��>�S�>��=��:��������5��=��>���w�=H����<�2���<�dƺ��\�AŚ��]�<�a�=I7+��ͪ>�EP>�h6>�d1>%�R>�����Dֽ5h���?K>�����<l�b��0n>��=K�1=Oq��ࢽ�����&\���]����=��Խ��m�I�C@���N�Ŗg��G���\\>�o�<v(>�&]�S���RO?ڴ,?�?�ƾ#�=gܜ���U?��\�e�*>�>�>�&=?��3�R>60��Y����=<�l��>�0��;��*�Yq��p�<도�۪>"=?�y^��p��ϲ<(�K��dl��6q��J?��>��Y?F.۾��5?f���p�V��_�=�fϿ�X�LL?����jo;NW�>���?�<#�1�>ͽ���Jg<��=>C�?�g?yK>�ާ?/W��%���>�W?|xy?�C?�n��E[<"�������H�>�螾Q��?v��>TX�>3HC>�$?F��$]3�]���@�?
���$��>���=�,?�"�=§ɾNv<��]�>���=kj,���ܾW��=�>� g־P���ɺ~�#yV�-Q���s?��o=(%>7[����Ǿ�ƾ�S>� ��y����<���"�?\7�?%��?�H�?P�R���F>�:�AG?�*2��Ap�ϕ?�V=�4����|�zK�>j��>��Ϳ��W��V��
�Z?�a�>��?<D?��?m�/?��$�t��N���)� �?(��=�j�>0�Q?���w�>�x����>Z.�����>̮�<gzg��?�����WC>�D?闌>��?߯n>�)��Z��.z��?k?�
�>�˾6҄>���pV����?�߿���B�kbe�tlH��4_?GSb<�~>W�k?b)?�D?v�
������>"�C>��>)�!?A�7���=>U��>M��������=��=C'f?"H�>��A?�>�����C��,׿E;?M�<�����$�[�5P?�>%?Q?:>?�;�]�>�#o�y�*?�葿66�⹛��W�5,�?�X�?��?��M�vQ?�!?���>��z����?d����b?�f?6�)�������=���|����><?���x<T�v��>�[@�wF��[��C?��̿N��/̿}��>{B���d�?�`���j?�9!�iiY?����>�B�>��O?V��?�t}�:a>2v�?��?�ߦ>��>o����>�d;���ɿV�Q?�]>9Қ=2�μ �>6���~23?�����?��>e��>4�?R�
���J�96���8@����)vP� �r�x?|,?FR�:�y�s�������ͿG&����
�����D�>�a�}^?/+���1?i���I��{�?�"#>��?���?۝?�M>���?H����J��B�>���?���>¼O>�o�>�������>:�����R�@��'�q��t�>�e">�$?7E�<�����_���?tO����?�C�Hg�>�%W>��"��>�w�t��>Q앾i(1>0N�ǚR?6O��6N=�0�پ���杧�>@�=2^>�47?w\8�^ *�D

>�P?%1K?d�?��[?g����@3�c�V�#,I?~���|w=?�[ľ`�*?+������,����!n��9#?���1��mx>�r�N���C�п�^��%=ʾ"!Ҿ6?ei1?�vl��K?��������>d��>���U��>�~����˾4T??��=�I�>��>�i>��OM�w�?y�z>��?g��>c��3��>R�>f����8?�$��[���|�>Q��?�NL������-#���c�P����p����?�>R*�>�>�!�>LK���Ѯ�.����^�����>�b?�;>\�)��/>�g<�+��_�=���s�d?�Wa?��=�@C?v��t�0�%~E?ȾqJ?�b'>+���v_��m��7\��*������� �+ ���h?�n)?~�����x>W���i�+�P�[?CAV�g�r?�x��?�a?n��>Ųj>Y�,8=�߸����?���>��>V���KGs?� ?�?}67�&d�QZ��7��:K���?ěl�v?,#?c��Y�A>vC�c�|�ܥq?���<%3�Η���\X�!��mE��狾\5�>Q��>���y�J�����#W=�
I<����n���-���=��?�����;��v�|�w��R��>d��=��N�Yѿ�8E�G�&>�8�����(}��\Yg?��?�ѽ��߾��w?�7˼�R?�(V?���U�w?��?N�	�?yY������8���F<��Y>��7�e�j=��>��>�?�y�=0|?z�N�
�,?)�D=#�?�+�=�U���X�?���{��=�=U���:����>�B���=(Q?��5?q巾����#�����=�%�?1?�U���{V?/4�Q�@N"?����t؍>��
�`b?g��%��eg�<X���l�C����;��B��ǡ>R@t?_�	>1P?4�?�X�>DP�����{�H���?]5/?��?�2�c��>���*���I?��?%��A�8?�t�ؽ��f`?��c��@8f#��S?G^^��;�?t�9�Z >���?Xz�?H�?zLW�(�?]U�?��p>FhL> ��e���u�b��X���V??,*��y�>��3?`������?Չ�=z྿ah��?$�a�H?E�>T�^>�.�iͷ;Ā$�N;�>r湽-V+>J�;n�>o衾����+,?U>��,}��G����>>Kw�=���1�c?��X;��Z?���=�ҽ�_	@�����1[?��>�Bh����d�>!��K�J�>�\�?){�?Qa�Y2?u�?�P�>�q�=ˈx�጑?�!�?=@{f�?��>���<�����p���<q��rξ���?�[�>��������>3n�?x���Yu�?20 ���?pG��0��`�`��y:��*P>�M�=釂?Ŧ�>˨�>`�*?�?�FԻu�@��>�(?ER$<�3�?p?�I�>�v�?4V�?��޾B�H>f�S>�_U�0�N>!���:�?���C��>�$*��?"� �2y���p��n+?�蘾w�˾�P����Ń�(V�� W>P3��'}> 'J��?��P>k�?��>�L��b���O�=���4�ھ�I?ĉ=ƻ?ƃؿ9:>xq�=9�k?Uܤ>��="�x<󀂿��>���=B�N��������L�q>���-�};
��hp?�ы>��?��C�Np?���l��=�J4?���v���:8?�V_?�NE�M|��ڣ�6A]?>I�?���j�M�a	=���?��>�F�>�s?��b��╿6��>&J�>:X�=u8�>����!��>�+H?�//�]��B��|�X>�/A�y��>��I�ʃf?��3�����K�=��̾k�>���eG.�#t�?lڦ�eR��jZ��ԡ���ĽO߽�'��ϲ��恔>�Rb�1�?�?�*��IU?�~�?�v�>�HE�	��aȱ=��=��?�k�=#7�>�	>.�þ�k?��<?��?U��?)�2�����~�>��=�A�=
�R��]�;�������~�f�.�>������>*�j��w��T>?O�X�|����?�(�)��>
� ?��[>�I>66ǾT� ������?�?͊�?�lپ�r? �@����un��0�=��������6 �
�̌پ���>���ؓ��u�?�w�>��<���?Yb�=���>����@�>n?l�a>i;�?���N����*?�Y
?&��?�l>��L��ѿǂ��c���y�]L3��Ҿ��3��8�>_�>Ҙv��翦%
����)�	�d�D>�G�?V�?s�쾢�0�Cts�T�%?�� >���>�<H����=��}?���S��?�(����>�'�p���پ�i�?�?{�w?��D?E��>���~��k��?X�>��]?ˑ���Sg=�Nо^�?�/C?m�=ҤD?ݜc�G(?9�X�D'>�??��̼���>z���]�>�Ƽ�RW>�,>��x���?��q?�4:��_�>3~����>��]�Vͤ?<n�?r0?���h4�?��3=_A��W�>�,=?��?( ¾1X��0lO?�v��I>���kh�d�;�-d|��3���Ծ�u`>�x�=
���!�ȿ�)	�uq��廑>P+w�����2�>|I?�B?�����=	�� ��V��2>����f�\?��N�M=�O�f�Ծ+�0��?�w�t�>��6?� {?3�<�I@�>��U?ă+?<(��[�=	V���>ڭ�>�۝��v��K >�A��8꽀_��=����>����jL?:!m��ؾ)y�>`?�����%�<��=y�'?�?h^e?��>qg7?����U��<8?��D�8ѣ>��=����y5���?Q)��K�`�����en�>P��o�X�Mr��#	`��ͫ�8���*u׿N燾,�?�>�?�/�?������-�M7��	">����m�>��
?8po�],?��>��9=K�d?>x���0��(6>4ʾE|�=�h��>����<�g>~@�&�
���j>ՖK����� �=v�Q���_�"�.��e���������M� �KJP>ݯt>�?>��F>�4n�,�������r���پ�����qR�u�9�fJv��_���1l���>f��!�]��V.��9Y=��?�9H?�Ej?!??��������ʊ2?��u?��a>�?w�����r>�Yd��/?�-�\.C���]�4���N?lOA��.�Mhj��2ȿ���,嫾��t<F�>���>ȼ�"C�?�U�?��>|�?D5�=ܑ`�1?�U>$��?�Y뾙��>�����=�XJ?��>c.�=�����e�=D1S��\�5Q����`��?T5�?�֩?�Q��V�>Ֆ�>��-?kQ�>�>o�$?VD>6a�>O#�~�"?',���?�|f�9M�;Y�g?�B����;�`,x��So>]��1e�6��Z6{�Hס���o�i�0ݲ��l�?�aҽ�3>�/�=ƞٽ��Q?�qH�e��?��7>7A=:Q�ؘ?@!�>�b?�e�?��ҽ$
Ŀ(xݾTXǿ��?��)����>,��={ڊ?����w�������/����ı?�ñ?��Y��?6���;x�?͒��I�E>bw�>��b?��+�z�8?��f?���?�\�>u�a?�	�>�G?�"M�����2B?�;�,�t>fe;?%⾫� ?��y>Ea3�s,Y�Z��>�m�p��?
��>�>��}���Q?�?&��>?�b��eH?�H�>��=�Ξ��QV��T��si��n��d��^�`�������~?97L>\��>��	�z�=r��=H�'>����Kj�>��!?��!=��^>,��#��>HB�=5?�̑>�d_�=z����?���}�>7�+=��8>��(�}B>�7��u����=?��/>�O�?~p/���>�IH>�:�>�Ҫ�Q�>�T�?ؕ>4��;E��>��>�c�>u�7�Hb=^���*�>'��dz~>h춾7�B>Yoɾ6���BW=���>iE���[�=��7?(y�>A�?DH?���>���>qW�Hp'��"��K��=u_7>3�)?�*˾-N�>�Sľ�� B+���!��w>l},��L��=�}>_���g�=�ھ�82����$"�o"=�=�> �<·=+>�x?v)������q�����FW���'��=se?��?��ƽYs�>C?u��>�o�>(��>X�>���d$�s�=��^�`v:��C'�o�?��q����w��0+������b����>Eq>.�,>������ߕ��}���m��@�b�m�����#�tH����Һ��l&���>��H��>��?�	?G�����?�2}?�)����辜�x>z=f��?m��?Bh�>����}�Z����=��?�&?E/������Vu����D?���>{u�jr��Ⱦ3�>�(�=C������m�P�6��>,�?`;?��;,^?r/?G�A?��i?� N?P+{>���?�
?�2?�ר����������<S>�[ͽ(�L?�EZ?jqq?7�>=Xھ5O徂眾D�'>�v�����V��@L��:���4��?�=����ȱ:���<��s>��\�����t6���>����z��Wd��I
?x?���D�=���>��-��= >�Ϻ>� �>��2��1�Aɾ3��>��|�5l�t9��w-4?C��>���>��>��I�j�>���F��>&Cp�?Р��=?�b?�����_>-�>?�Y�=`��=H�$?��y>��>�i�>���=ټ�=J
/?�f�>kb?�<f?Jd(?t0>+��?\*?z�?L��=��%�G�¾�S�n+@�6?�@�侘hr>��ج��\�E?�S?G�&?��T��μ(d�]��>�ME�;@}�����d>q?LU>���.?s�	?�j�>(W�>�c?sW7��`Q?�d{?��	?�Y�?��]?	yE?�h����^�O��i�ݾ1k? p�=塬<G��j���U�>��6�~A�S�|�޾��>�Tg���+�B��%R?�2�?�(����>���F�?.���פ���"S�e"L?��<��徾�Eg>qy?l����G?^�~>&�[<�����0.?ZJ�>�l=4>����5<Xɠ=�ݾy�&��8���(����T��>�O���'>cdA?�2><�C>=�?-�A?'?W^�?O��=�	�>q�d�ƾ��aY��R��8;�>��{=�S�?1�6���?ni�>����7>�?�I>C�?�'1��f����=�`>�׌��Q>�:˾i�?A4�)��?c�p?_!?ǌ)?��?T?�Z?sG�>�#?RN�>�0?P�6?K��,/?��>1��>����{
y?p�>��>`��_�F?�~?���>:���d����>Q��=|�e�%�=>U�W=,ի�S�>��U?�5�>�MW>��,>�h:?ې�>��>�Tؽ��>�a�> U#>�Z�?���>	��?�������ve��뉽�}?�+a>�����T�v þ�	G�>; ?�߿;ҍ������I�p��>�+����s�'�/��΋��ɯ����U�ÿ�5^>iي�� �?h��>�.h>L�)?O<?�Hd����>�Um��;>e�`>�b�������?I�sk���ڲ��D��/�&�����H�%�Y��=���?���$w��7��=�<��ꕭ>��=2��>y����L��U��fK?"@��+@�ķ������h@��K?�Z�?<���[?�o?m��>�1��ƅC?�b>DBA?>��T��=ź?v,?��L���]��>
����>;��>�~N�[Q]���������M��=��>&���}�>�[�>&bG�|��?�_?�z>�y�7��>���>-[+=L;E���[?�AL?G��B� �	����Y���c�>�L�_?*?Bf%?�_>�*ݾke~?Q�~?Ձ�>��|Q�?Ld�?䥠>�z����Ӿ���>��m�jG�۵�>#T~���I?�>��=����9��e�T�q>Kf�d�����4?m4>������>V#Y�]:>�ފ�z �>\��=
dc>�j@�bϦ�rL_������t_�Ǹ�݋�>/�?������>��Z���?@>�a�?��>�>}B<����?,^�>){�?k�l����	��b�4�L�j���+D�u������?�ވ?K+x?`�+>=r_�X��>��:���>����G/>?.:��	.�=�羗x��3�]���u��	�7����=
�c��蒾���>}T,>���>���>�Au>i����#?@�`?q�7?��?b���ܿ8���3�����(?d&Ӿ��Ҿ�?}�E�8?�������������>>�����&�>,ݽ��:C
���̾��վ�Rd?�W�>E�����^�>ԟ���*�=x��pQe�+C?�[�>�R��1V[�K�?|��>���<��>�wR>
7.>Ϗ�>Cɚ��>O'�w��҇3��^O?�^�>?e?���>�)Q?��;�8Sм�-ᾨy���)�>H��O��)�t�S�r?�y
>˘�>X�(?�\�?��?�Y�> �(Ӈ������^?����W�n�7���??�f�SP��q���8�>VϪ�5d	�z��J?)OF����t����M?n�e�h�M���1��˙?ٸ�>B}�&W𾟌�=Â�?��>4!A?@?���=�S�>U9&?�k3>?��aI�>�w���A��\@.��>.{�=*A?D��>�s>&�]�>g�۾���=_6�>-�?cX�2(�����w��]C����=y�|>�Q�9v�<A�P?�1�>�n~�yb侾���qz?�%c����=���k�?{$�>��=>�6< ;j?�M����>{��>��F?�2�?��=\��>�ýCH������q�S��@Ç>�y���]>�JR?��->��(>��ο�5���e����?��q<�ǘ??�������۾.�Z=��!?d��p?��>��<?�p
?a��>�#@hzI>����wzĿ��-�H�>��:��X��z�>�E>"��>�>�sf>ı�>O`>�MH����?���N�=��U��7���d���H�=j-?��w?~��>��>�>P&>���>?Jů��� ?�O/����~l��.���t��a?�l�*h>�*�L�`>����⽔?�.��"��>B��=�2/=|�1?��>�J�6;'�>�������>���?��Q>�3��xe����ٲ?| �?27��J:D>j$���l�/=䝚?�+�����Q�����k�)&@#�?�O?!4�>��V�ˑc?�S�>�*ľ��Q?���2	��J_�=���>�"��?�Aξ���>G��F��=�?-�,��f?6��=&sO������0�̓�h�?��G�q,K>�a�<*n=�3׽c�?�"!>�D.?���
&e���>�? 큾[�_��)�??�t�>bze�����2�����>LB��]��?(�?���ʼ�CpX�z}@���'?��H�?� �>��>]G#>r>�z�� �?o�L�J�^?�1�΄�� n�>�=
>ぢ>�[�<��u>�#w��)Q����>ܜ*>�z�ia>�	��2���<گ>W9^��*�U<�w��?osY?�T{�L*����?���� ?�U��%7�?B����]<�m�>��?f��=\\�>}Ё��?�<?����b;/���=oV?;��>pl�)��>0����>�?��*R?z�a�x�����?)[#?AZ־�/��A%?LO��Zg>͹�� �k?�}�d�U�
B��&ϼ�6->��	?�g�ϝ�H)�D��>���=*p'��\�?�ׁ��|1��B�~e�?�Qھ�;b�>�*7?�"?mA�?��|��[�9:�˾����E��>6��=k�&?Oc���־��b�}� ����f?�C?�����P+?,K>���>��?�L���?�->c&�a�6���F>0��_2�>�l��鰾�t ?nD�>��)?�
�<TM�?=���	�ŽI?�K,�?�5O��/�>����b~�?3S>�I�ʹ����?�ح?e��?�i�?Y�?a�r��GO��ց�
��>�ݒ>{���y��#C�?�/U?ܼ?Q,?�Ԅ?��$?�_�>͎}��C��󿏪�>����>���>�-0?��3>�u�><��?�>↼?�h>V�S��,ѿ�y]�	*�?�1�Ȼ�=p�=�1!?NU����?��ý�w+?�8�?�~+>'~�KX��ʍ�>�ٓ��d?�	i?���?_�=�[;?|8���>��_�]�Y��̾㓞=f�*���<0���H��0z���?RyӾv����d�>LG���G���.�uꟿB�4�6V��\�=	�?V�E?CK��Q�I�^`�?�\?lD}?�gG>@)b?���>����$����}>^#�>fX�>�c=�`f>�6u9�]E?u�B=�ׁ>8�H��?��f����>�ۃ?�;>�������>��?�㑾�L�=��>�<B�u>�!Y>�D�ص�=��I>d93����>�u�?�@���? {@�4F���W�+�>�@5�p��?
"�?~�8������>��䀃��9>`aP>7U⾳N���<�3�$]���\>:�>ヽnھG�>�ͅ?/L�>s����9�jҧ�J!�D8��¾��Ӿ��E>�������=��4?T��>��=l���۱==�?� ������u��>��G�F"žgξ���=�(�?~ �\A(?�Y?�Z[�ݲ>���?�9��-s�>��Z�`���i<=gu?�8d?�E�>��F�4K��<�
��Op���G����=�s[>��
�!�|�^��\?�<<@!?���?��?�/�>)=?]8��%I��`��~p�yrk��y�=�>�O^�?��> �?,&����gK�t-?������>o��>���> ��l��,��=ջ6>a׾���>�=sP�j�ξ.�$��ܽ�?�E��<�?ig?@l8>��?
�
��"����Z>�;�9�D�:��=��?���>9�>3f��Sž�g'?�`g�G֢?]¾�]��?�\r��J�M�4%����?���>�>>��O���?:����D?X#��J�?ʎ��w����8�wT�?D.�S��>�c?E	�����jn?�f�>< ����P�0?�#�<M�>�_�A>��	�H�N���Z�c=�A=o|.� A8?��?ԥ�<������>������/�����y���i�^q<�q6Ӿm,?������>�#k�..?WT�?�ݫ?:��|-?Os �5+�?^�G�4�)?��F��{�?G���Q>_Rb���,G����<=��>�)9?��B���?���>7¾��3�C?=?�7��w�[<ʾ� +��[?����G#>�Й��_E?�_>��/>�����Z?�v&���E���"�*�?"ᔾ���?�����>�E�>��ɾ�{H?
�?,g�?��%>�^3?���?VC�?��?8F_?�,D?� ?Ś?�$��b��E�l?E�?̄=�ƴ?�}?d򶿲�����?K�u?@%"��HC�۷ﾂؿ
�TE%�R澝����P?n[X�?˸>��>	��>����}J������Χ=�?��>��%��d�>m����\���3>��1�=�U!�v����;=ל����?�+�����=:�=���_k�>1ڈ>��?Kg?��?������k�+Q�>f��9�>�^�?��>;�=?�̽�$���=TE�=,0,��*���?dɬ=N<�?{�w���ǔ-?�/��n8���Ȋ��y?�� �$I7��.�?2:��+��N?��|?�z��L�/??X��=������+?�@	>���&d�v����?+`?p,�?�޾�a�/c&�$�?�j?(��9�㽉�?��[?ʃ��
?)5�?r�ӿqsP�`3y>`$W�U#>�o�>���?YA@�!.�Q��>�ֻ���>�7�>:ḾB��?=��:�cݿ��>t"?�^ܾ��"ϣ>AS���a?jE]��b�>���=G}5��o�?��ԽP��*���e�.��?��z?��	?�~����W,f���@dŒ?G�u>�������Ϟ>�������,��"S> !�?��4���{>�����׾JZM>b!>�<�3����D��$?.�?��!E��N�>iڻ?ofܾ<��7��/h4?w[l��O��>�H������aS�k
���̾�{�?�Uy?�P���>%��<(�t��0.�J��Nd�O�l�����*Ҿꕡ��W/??q�? �elQ?O<�BO�?�l?l�>�c`?뤉�����#w:��`̿� ��>�>nV�>HU�y񒾎�?ش˾ �j�?��>kN�>�ǽ!�8�[���@��>��9��uϾ
�i?1�?���>L�=*�?�A���6��.�,1�>�����?m�6�v�+��Z��t�_:���]��0z�y�{?���d"?��0>Zm�>�	�>���>����*h�t�n>�FH��]WU>�c�=�eW����=P�J?R�M?���>W�a���q�[��GF�:������?�!��t�'��j @� �U�����>���>�*?�/�>�ܚ�q��>���? �d��?��>�JԿU8.�5Ѐ?s煾:N��\G�����?��8 ���K�����?4�N<,˦�u$�>0�=?/���wu�?�H>([�?1����:V˾���?���?[.��_?�H�>]���=ou�<�Ø�b�>�6�5ĺ?�c_?ML?�*Ծ)�?a��?�A�i��D�>�u?Sjh?]e�?��z>�:�?� ?)>>{�->�-�=k�+�kϾ<���>��?��>����?��������j���?����� ?EVI�X9K?�޸>�*R?d4>��?���q���DZ?!)���>ټ?R]	�ֲ����ҿ,b����>hu�>_>��P>�D=-���A(2��Ծ�	\���ƿE��?��_>-��?��Ž.��?�wg>���uSj����>���?Z U�S��?�q]?���=�D?Z���s�,��l��Yu���m��<5��)'�?)�>M�Q�}�P���Y�n�;E���d��j�
<��a?+��<�н��>| ?Z/e�Dը��<?�J���m�?ӻC?6�_>��H?� l�Ur?|)=��>,r.��Ǭ�A��V�6��w���\���[Y?���>(�`����cH�� �vTм버�k����J�{��#?g�@zc����u���n�L�Z�����$k�>��w��,B>骼?v�V?ߏ��!�?9`޾Ze�=�ػ=�Z�N>��1?+Z�{0�?�!N?��?r�>���?��������wV�>B����?j�>l��>�?+�����?�;N=M!9?0>>�R�;1�Y?�=�!�0�>���>OXO?~�=�Rl��S?���?0�(?��>��Z?:>Ҿ7���;?:2���#v�Iǈ�}%����8s�� >������?��=������>X��?Iؤ�4j>��+?��>��E��W��^r�LHJ�R�?U@l??F�?%��}��>�����2��M=�/ ����>΀>��<\%�=@۞>s��>X�O>+�>��T> ��>訧> �>��>��>�hD>���H�W���?׈ڿ~#*��X=@q���zq0<�T־�T@����x�><�n�?���{й?�����?*�=7?5��>8�%?��
={���.���×?5�i?ǿ�3̾�UK?�?:�>�� ����=��!��O�?;�>؁
=���pW"�þ�J��
QӾ�>��jx������/�"�y�����X��H�XaӾ���9?���d?M�?2�?�E���}X?��_>/g��ע=ש(?�Z�>w3 ?\.�?Ga)?��L?4jh>���?pї?�/��)
��h2�?#����J�=���]6?�FY����=�u?��Y?���?�i�`-��(?8�-?'J?7�
���z=���?ze?�t��*?�O��<�ߓ?8���
?��ż��?��K�?�[4��l��-�0�R?R���� ��3�._@?�����p?�Oq�<�E?tg�?�r?��?y{�?�7m�?Ȃ�`bſKLR���@;��`�+��=Оڽ(���_ԏ<J3�L�?��R?��ӿx���V���?Qǁ���k��3g��y�?��X���>(��`� �N��������Q����>*���k�>lh�=Ҹa?7 Y��rr>y�z>�w ���?(�3?`�#>*����,��T��Z�r??ߜ�u2?La����>+�r���?A�>?�K��>�=��R?R� ��1�<��=;���4��j��WR(�����|&�HT���[�<_��>�o�>+�F? )��wœ����>��你�b�%>������?���?1sʾޚ�>-B�>�%U?+&�>nEM��E2?�ٕ>]|>w�=�+>��?��O?]�@?o?	��eA?8?ّ��{fV�D�l��"?����C�;?��)?��U�TE ��Q^?�7���0�>rJ?�\?��n0���>�2$?��=?fKe����?�J�>G�B��>l?%Uz� )E�����0����=�dX?a!;�oV�/ߝ>�f����?�)q>9޾F?�]=>��g��9�>܏��nF�<Ut>ͥ�>���>̕�8�>���>p^��9e��>܎�c޺�f�h�y���!=<4(?�i?#=�>{�?5
>�����>���?}�Ŀ��(�D�	˄�����ҵ��R�;��H?w`= �]�7F�>�ԑ��T����2�ޏž���!��,w�?:[���)��H��yȽz�3>�8.�+V&�%΍�h+A����?d?��r?׾�=��ݾ7�?�=`.&>PH�=/,��
���Ȳ?i�.���*��'\��t � �G?G ��D����?C��?K� �)!��#<��>ә�?ȫ�>������;�>��i��x>Y��R��{0�sQ>��4��l���jg<���W�?G�>	��0�*�Ӝ�?�)�>�
�>:�t?�	��-�PP2�0`9�h:����)?m�>�q׾[�>
��*�y=]qJ?{FI���h���%��eҾ؉?e���U~ �A�?7t�>Os����ַ?m)��c�+�i0����g?�n$�4w�>����K_?$�����?d�{>�B��y��է?_�?��>������=�?�A�>�����ľ��B����>�����=jT����ſ�1޾��?��?��ɽ�q�]_����%?e�>z�q�ɲ��*��+^��2���I?�=@A�z����?(u�?]�>��z>�N9?�7�>Qt�?�w�R��>�+��UQ~?��X���Ͼ�g��j(�=��C�@��>����<?��>�Y0?b�j?x�*�����pK?dQ?���>�*=&�����?�!-�$H]�Ѓ�\�����4?�,��^Ͽ�n$�B6�?��Pѿ:y(��?^lV�M�_����>*��<;UA���8���?�k�?�-D?�7y?r�]?�Z?n_�=�p�>D�\>�_?Z���h�?���T.̽)�5��?����?�2>��?j-?f���g8?�C.�*�?h[�><�Ľ�2�e劾 �3�{�?Ҹ?��m?/?)�H��a?nVG�|�>]4�=��)�Gb?y�o>5��>% ?e�0���%?}��V�]��h��T��ҽ�����z@��KϾ�;�?l� ��>8콾}�r��:��s?�?CA�?�u��)B�h�y?�� ?�=<�*?R >�4�(W?��2>�.�<�ֽ�r{<9S��O�?X����<l?�,��^�?�Ҡ?����ο\h�=�X
@.�}>I�这�@?���?�����?�W�?!������>ǠP�H�>���>9��=I���l?^�`���>#,?���> �u��>`-��)/�?K�?��\�@�{�?g;�?�� �lX5��S����?�0>������)?6��?�0�<�J?md�?S�=ݪ�4�.?b����{>��K?q�h>��Q���#�:�>�CX?݀���Y�U�����J�;��WN?4<>~S�-�9=O.->)T<�#�>>��?4"o��d������]�v?-��?����i������u>�fa?�m?�FA��-��a¾��j��X��I�`?g��>�?�#���ÿzݹ�8~�>�O?[�>������?#�g?p?�ㆿG]x?��=y�?P���ھ�(C�#/l���g�x'j�.8:?>�K��h:7f0?<�?�ԍ?�tf?1�_?X�0>žA�ڒU>�/�w�!?�[?H�'��}��%�S?~T�>�p��?/�?I+�?�l,����>8��.�?(=]�e�>�s���|>�t־q�#��r��Ue�x^(��r��q]�?��D?Tt�>q���A+���\����Q�=m��l&I?_�E����<8��>~��>yKV��=ſ�ר>��¾4U�>F�>�7�=/t?��q�P�!�i��'��=��ϽX��>�p#?��g<b�q?]˵�j��>J?��-?Id?�풾���=x�>�=z��%?y�>셾��>�p�?!Ǿ � =�@�1&�>C��=hx�>&(��&x"�y�1�I�S�1��>��E?0|�>�L��^z���)�<��"��Ft;�z�>�3�?\��?�EG>d�>M��A�۾_�M?*�9���E>6���7?]z����S?1�����?L�O�1�\�p��>�,�??����䯿U�½�{@L�=��R�Ĕ�>ٱ��m�?r�= ����h��6��ނ���?�Y��蓥<q�?�u������4?,�_�tq ?�r'��@>}��>b�%?�V�?���?C�w?�(�?$'�>��v�T�O?(��>}ֆ>��=�q>�t�>���L޾��>">䎫������/��(�8C9�39��'��>��f�KL>2x,>��G?��>�H���ֽm��>;�ƾkz���O�r�)>L㦾�By=<�>�L?N $>�k>�|7?Q�<����4=�P�=Afn<\Kh>n���{���	@��_����0�����P�=�*u��(�=Ek�g�Z?�FC>��><�v�Wǽ��5?�a�q�c����[�����Ϛ�n�I��]?	]�3H�j�/Σ�Y�>2x�=�m)>Pp?��O)���M����2�\%5�0��>�>���>!� ?w:�?<�??g2H���o�����c	���2��q+���r��?�?��r�ɜ��,!?�ޛ�*|�
Wp�M�ᾷ�n>ʼ?�����>���^��?����h܀���>���#\�>�R�=k�7���,?&x�����n��?.��>s)��.�n�|��?a���%C?idi�Pș���>#�?��>��?�-�?R �>����	\�>.����!
�>�A^���f=��>_�?�!�̗`�`$p?ПѾ�D�'?��> �>e�>h�F�(��AV���Xq��l�T�e�ാ5����~=-Y�A>��?���xQ�>�>o�g�'vA�y�?��e?6�Ⱦ >@�4
��?Tr�2?���>�+"> k�>��L�&me=�5Y�3��=����k�j�;��>��>}_�?[�>�ڇ��緾�	�=��}?Y�I?l�n?�׮����=e!R���\޾=��>?6ƚ>�.�>�x�>멾V�s��.��?k�=`��E#?.��>P0��:R��U�?>Q��>9cZ>���|h�>\e���C�2�>b�;?*-����g<H�>��һ�*��,?��O?i��>N���8D�>�>W>_����ѽ!� ��A���2�=�y����龈�w<�=�fs��Uh?�j�j�=�
�.�m?�u>!�="ܩ�3+N>��K?��>��Z>{��?Pԅ?�z�/(˾Aw����6��66�+l��~�`����>�aI��Ď����lǾ18Ͼ쓽�a>��=�^p>�r�=x��>.��>��n?�?���Q2��	!?��2> 3�>� �<U�����|~B>|3ӿ]6>�kc�)�K��LI<s]>u��]?H8p?�ݰ=U4>�.���%?\m�?��C�_�I>`1�?DOA>s̚?��>��{>_.?��s�D_��{p��>�e
��C���{���˭�<��tþ(%�>�焾}9����7<@>ͻ�>ؐ?t5?�6?xҜ?]�>�෼Y��=f���J~���I��"	?�\?�7��V��$s����M�>���
�>0@�>f���=��W��4���+>Z������L>�[?[U�\e�_y���R����>lj(��^оT�!��B�>oOM�h[�==�]�5�b>��5���.��
{=��]���Y>��>w�>��������<����
��N��*>CD㾭�&?ؾ	d������� ��Z��=���>�r��B!�RX=>X�?AU������"���ٽ�k%��*:��W7�ku��Ǽ?v�?�?�݊>'�>�ɍ?X�n�)��A�>��K����>��T?���=�E`����>#����SE�/�S�e�5�
�R�8�<�zK�dfn����=�ܘ��)��oO��8N)�-Q'�ľ��G�?�y�������"��$ֽ�,&��._�9i=+d��&-����>�S8?�w��l+���E�S�/;����V��n��j线��������D?;`���>��>¤?8&F�O��>���>`�I����>~��1�NŽ��1R�>V�?]�=�����p���j=py�"ʃ�9Ȯ��]>bd��_��x-��a >׼�\m���->?>�H���?%�̀D=i�>�.I�Yfq�MC�<�>��4���c��S���>���Mt�R�= ��=Zľ���>8T��"f9�(�9�*�?�g�)>&&�U�=��>��ؼ��?]�"�$N	�c6��<�=�ƾ�U,>_��h��5lǾ݇�����d>�}�=�Ua>��?F"��G����=�6S>H���^�? ��>�Q�H�@?܏x�H">�ax>�$D?C�;?S^o?��[?2��<�s�>G�v��$?�Դ�*�h����	�?�}��J���	�>,�4��V��]�ɾZ�c��,�?�;q?I/?�d�?D��>;-f���(�hC�/�X����&7�*�����Z��ᅾҝ$��¾Ev������>M��L��ά=�����Wh��O��[��>fᎾ~�K�a�f���> p��O=�~�����X�*��=�RL��]"?��?�м�'5=Sr�?�"H�W5?7����l�?�(c���Ҿ��?�o��#��=N�/��痾�&#?@��>�8�>�FQ?��>��Z�nl���]�>�>Y[��TZ�?tQ&�b׾g��A���4L��a��=݀>��?�3�>
Sｃ��>\@~=[�\�/��2��>���Y_�>X"!>�}�����>ՙ\��o>DU�>��Ⱦ����	?]%I?�S�>3�+��j?z�t?�B?��58�B��>*�?��i?L魽��J�Q��>l��<?�=MC�s��9�3?6Q(��*���`s>c�_?��M?�-�����=c;q�$�)���3>Q۹<f89�/��=6�V?@#>Z����X+>�H�?[�>��P�3$b�Z��ٚX<̿ʾ�L1?�Fξg?�6��1�>���>�3>���?�@���J	>�D?7�W��no�q��=��?� ?��ɽ}��=.r-��=�i��>k<����50<|%�=١���>�@��
��>�+<�	,>�bо��2?�f��Ȍ��`��~/�B�V���6=���=���tӀ?>:A?ci0�B+����J��G8�	�>
D��S�S�T�����>WEo�Cn7>��2?�[5?�o>|��>�＾���>� 
?C�2?;��>���>�Y��?Wؾqb?��P>�
��w)6�gB�?.ݓ>3���h>	W@�� ?����2?V��ۧ���U���<'��
?L!���߻��ľc:��$ҽ���?�y�>�M��{�a>��߽}��� -�>�Ȉ;�^P=��>�rۼ`�?��z<�?5P>�&?:�>�d���f>Թ=�a-�z�>�	��M?�5X�ݹ6?j>�ξ ;�>ԇ�?칾��="�� ���h������0>=�=��<�1�Ӿ�T�=��ʾd>��q>�[.>�|���#>��!�=�:?s�ֽ0��>;B�?��&���s?6��>�����C>��1�&3%�I=���$<�\?����A>7st����>�d�>�S1?�E�	qE?;F�>1\�� ���osx?�/O?��E>�v��f(?,�y>�u
�|Q���7�kؾZt�yힿ����T>v��>
��\
D?M�?$̢>�\�><	?B?�,?��W�d�����>߰�?��>3�>��?�㻾�}m�(؋?o�U?y��x�?��F>Z��>��Խ�@=��A?��?�* ?�"?����¾Ю:��qd=�'���Ix��T�>�J>ǣ�8۾����Yk�>��ʾ۴��n��ޘ'�E�>h�����c>�0�>�1v��7�>5OL?�;R����>W�"���O��s輻���$�0�r����饿� �PV�;ܐu<FN�>s��>Qύ>^]d?7�?ͫ
>.4�>�2�>~�?_�����?E�?����ȳ��w��������rӰ�Nb?nO��gr˾��t�=cy�,i?�RL?���� ?<�����E��@?�+'=�kZ?��?QH??�4>Cڻ�@7?[��>�7?�<V܂����?�]�#"�?���>(=?��>H�m�JU8�4��=�!��Ԙ��R>�,.?̃M�]���{J���v?��<�O'z?�a@?A{��_ލ>����y/��R=�,&�#f��f?M�ξ9����� ��`�@?E�?��?���=yn�>e*9?9�Z?&N?�}�>y����<��G?�~?�Q?"�D?��-?������TZ�p����ғ>�4	?�&1�an�>�)��W\���.���&?�=��Z۞��&8�\PK?�@?\�?pU�?H`�?*��݄ɾ��>���� ����>��|?NS���i?LT-@s=�?2}Ӿ�4���>���=����0�g��^����;>��þrJ���'m���>���?�����پ�i <����k'�>��}�'�?��a?��3?�#>(�=�?m?4�=��t����>�{���^Ӿr�>�C�����5ȾD%��˄>Y�}���Q�Ч?�<p��&���J��f\?tZV�����g5�nY���<�LI�?�7�?�w�?��?�6?>��7����d0�>�Xﾤ�=id����:?LU��.˺��p���>�L6��|�rE���i=��o>,G�>׊�>�� >�\;?�J?U��i7�ҶR?�4ྗ/>��7�:�n?�ᔿͶ�Ug����g�	�?HR�@Pi��C ?J�>ς�=M?y�P?��@��\�i�p�n?i@��@�A$?������>)a?��߾��?!�=8���UB��63��"� �[�>����s�����I�?�����<^M�F5����������*>!�d?z)�=�$�\<��O�"�ƿ��d���r?��@{'�?�#?��,�=X�>U+�=yϨ>���>�T>���<����ﮫ?x�B?c?<I��p�>GcJ�P��i�?��>�����\?���:s<Z�ѾE2��"f��ws���>�3>��?0>�2?����b����?1B?v0�>嶻?�y�?�Ј=�m:=A���g�?B�����þH+>)�'?[c�=>^~�t�{���3?�繿y��=x??>���u[M?�J&���_?_�����>A�'���z?ngj�9�O��w�#�?|��>��<���<^?;K?񙆿%�??	S?OT�>+�H?8�>���?ҽ?I��;@�п�y�����琾̜
>T��;q5��J�D=?��?�t7?��,���6?��?�V�?����仾༇��!��)v�
�վ&�k�V-Y>�k�Yy���پZ�>��>?��=��=���
#?����^^�$s��t�;>;�����%��O�?�Y�>��_>k�>}�>��V?ne>g�)>�	>�;1��Ij��k��^w�o����&>?T�@｟냾i�Y?q��?��f���>=�2�o&}>3������?=�xx?�X��}T���9�>	��>:-��J"��0���C?�� ��'���~k�H�>�'��젿@���a�>�]>N�7?6��?�C?���=�Z<2=f�?������G�I?9� �fvd=�'��6?h��>��J?+�>�����l|���5� �D�Ŗ��<� ���$�U����m���[?E�>y�����=&ĉ>z*�<���>B�>�ΰ�|�A�����?½��<XJ�
�M>1�žEz?��k?���^ܪ�-��۷�f%��������ܿ�̷�en?(X�>Kr?�H?+�'�|>i��'�f>�p�\m��|�F����>sB��z �%�*�Et����`>�?����F�(�:#�>��V�!�A�0�����ʾx1?�K�?�N ?u%>#�c?��'���?!�T��ǅ�p�n?�m=�|�>�(ݿ�y4���N������>���!i��&׾��=Y5�	�Q��{��p5�=�u�������?mu�?��սW�8�m\>��e< ��>��>��s=l�
?�+=%�8?���U�>�#@L��?JQο�hs��̇�v�տ����D4��^b><�>�$���Pp?x��?^�>{&�?m��ζ�?y��?ǟ�>!<X<���� ⁿ�	?�H>��~�P��<������ټ>���uj�Ŀ4��fa=4�⽙	�a�Ծ(��v">�K	��j����?���7о��j�(�9�����Ͼ!�W�D*��;\��g
۾0l��H����92?1%��Y��:N��8���ʡl��􆿸+ѿW7�W�ϼ�7$?A�Y��xҾ|<��1��[F?���>�_ӽ8<�>���O��>�u�>=�?�?"??j)>)ٻ>���?�13?��7������i�|���U��>�Rپ�@�?͛>ڒ���?œ�;P,?�A!�l�?�na>���?�B�j��>5G�?���?CvS�f.y�n��>&z
�(5~?P��>�*�>q{�Lx<?��8?���?пe�|=��j?�	B@��@��?Q�>���=������|���L��8��ÿ�Ra�ȨD�����c�(�?_�<#��=-��6�&? ў�� ?@�J?���=�q4?N�>'�?��V�X��>:���7jB?Q�����䂿��?o�&���8��h?]�U=כ�s
�>�?/�?v����a���|?Ƒ@�����j�>��)�������>q��>Zd�>�q�>�/�3wL=��>5˝>yaվ{MV?�� @U��?�JF�;�
q���ȿ��?�CR���?��$�F�?��n?��?�ha��,����>i��?B^Z������+�=�P��"��[��z>L=L웾6Za���?x��>~�w?9	�>�?��>����R6F?�:o�v�a?���(G@�c-?��̾{�?)A��R�[?��+?q�|?^+տ���>#�x>��qƿ�YL��>�=�b}>|���l����r�Qb.��+>W�<rc�>Z����>�~�>�wq>���<Yҽ���>�)�\�|l�<_���5L?&��A#G�k\H>�=S?r��?0����[?���?7�#?�])��\�ă��[>\K�=��� �B�)�p�X�=����=Q,���?�^9?�-�;v��������?1ح>�R>-�?�6�>��?�!g��R���ل=�F?�^<?6[�J�>m)�>�k�?��c��w����#>6a�ɫ;�D~����?��7>����M�?c��>���>�U���>��Z?�N]?[����Rc?*@!@� @ �-�˺>�%��>3�A?Q�.����Ɓ?g�<>���qYc?�G3?�A�?�rͿ�ꋽv(�0s	@2>T�L�n>�^l�IH ����>�F>���I�%?��u>�󴽽��Х��m�?%��?���?2}?�3?g4}>�F=ux�>�y.��>�܈?U�1?�p'��XʾK,ݼ�%@��>��y�=��H��V>1�Q���Y��N;��ZQ>� ��bq>�q?D��?9���_��>J�#�2D���eԾ���C�մ@���?��@�>� ��Rþ��־�if?�I�>�Yξ勵yq�>y��?��>I��\;��zρ?)�V?Wj���0��Y>lm�>T�����:���=��?>2��?9j��|ֿ^�
%ν�m�?� �?7C��T*�:dK?75R�ˆI?$�>`*;?i�����O��6�?缧?E�y����Z x��+o������.M�>q}>���<������8�&��$c�?X$>E�=�[��>��:�-x轈Þ��岾�"?I��I�?zΌ?P�>��
=8�>3��i�������ͼ�����d�n��ԥ�?̨�?���?��?8y?��?�����?x�?Ζc>0�#�P����>�
<�bn��(~�=��>���8�����g�2�1�E>ɻ��o��=NN?�:<`|2���1�s�b���R%h�n��<)��~ʚ��J��6g[����f=Ⱦ���>�g��?X5�=��>�?�>����?0�<��>���>c!6?�"J?(��>|����K��<�F�þ@�iW�����Ǚ�>�;?�KB����??n�[?�8�e�?\Gb?@�h=���>���>���=�6�>��w?/U�;YW>8�y�-�??��� 2�=H-���|�>�ô�Y�>�]�X�8�?��>(�E�B�t4?�6o>A�$��Q�P*=?Tv��R����� @g�?��p���IP�<T ��Q����ʘ�gӐ�68��x�T>����	n��٩U�Ĥ�K�=X̾9���S����ޏ�>o�h?�[8?F��>A�1?�zP�Xđ�`;>��*?{��?�g�?� �?�7����=[O?�4	?Q?�]4��nټ_?�F>f�$>Ķ�=`6�?�C�ɦ��o��?�T>�V6?��trQ?)�Y?��>HȔ>�&�>LI7���?��d�Ⱦ^��gy.?��D����>���=i�{�Nq@��7���'�e����=��p�D_�*���h��=��!?�?r�>l�T?N�?�7���nR?f�?�:L��̄?D �=�<&��©���>cE�¿��;]G��ö��	j��b^�ҍ4>Z�4>ܾ��e>��>����*�r�wr��\����7>g�>�" ?��z>�A>[��y�c?�
?^b�>C��>*L��]䦿��G�7�/>��D�Ԉ/�@�d�u�R%�Y׵��	�>l8�R��#l���>�&l�y�?��>|��>Y�Ͻ/'�>$�ھU$<�C ���O�.<1�����7N�rώ<�QC?�|��dF�S��t����<��l�>��(����>�n�=b�=Z5��i.?(�$�f>���$ >����U�u�n�)����>S?��x�s@=rO¾���<�΁>�4??MYp���=��E>@Ͳ�p$?ꦶ>��U��>u2?1�>����^،�o]A��S���>�&H>��>֗���w=Ƃ?~��=kQ��T�=3 �>��辿�V�������>���/t<$C�H�>�*�>_=����ma���y>���M���'���������Y�n*��G����>Ϯ�=��=Y�l���>�i���;��#�ٽ�Z�>���=�����?D)?n��>;
�>�N��>�����S�U$A��'�>p��>�� ���7��q�>�X��>�����IT˿���?�&�g��C�>�\�?�u�a6��?T@?��_�i�
��G��NMp?��+?C�/?Zs�=�>����xDc>{�y�z`&�*9���w)?��>�@ɾ�hJ?��?u�&?���>-a������>?kM�?&;3?�x-���!> �=X�4�Gv�:�C��=�#��<�y����B��t��Xz�(�3>��=�)ݾ��r�G5����@?���>��v�V�0?٫?�qS=�aI?�m>cЂ�Bqz?��>�%�!�9���y?ɣ3?�h���o��؞�>\�N>U]��[�Ⱦ��_�o�4��R8���]�81�>�tp��wc����>W|�>���=������>ΜK?L�8���`�*\J��h�.��>�y>��=����}Y =柿+!>������lݻ��H���X�0�.�X#	=���>!ɰ=��n�|�=�3�>7?o&�?o0�>u�>*���[�>^qսڝ3��9o���ս�����R`N�6o�>\���Ϻ>�Ь>�AN��j���m�>�G<G�~���f���a��>l� �m��kt?8���wD�>z�����>Ϳ>Z�}?��=��!���I9��������?��$?��߾���:jY��]�>��N>1a�>���>ì��ҋ���U?���>�x��_{����&>�U?��?X�G�Mp;�n�f��u?q3�> -�>^d8?@c���zT�CI���M�6:ʽ�.���>mg�>���>�kԽ�7��<g�ך����XX>D�>��?�w�?b�q?EA�>��~?�M�>��>��1�fB�>x�׾��ҽp�%��>R�Ⱦ�^g>��>i~�^��>�i�:u��<Ł��=�1V	�W5�m��/n־�&��Ɂ������\���#\��gJ}�]>j?�#�?�:o?9w�=W�?���>"m�����_w>
)�R?۲)?��l��~���ǵ�,^��2�X��>* ?!�?4?��m?�q��$��<��?�Μ>lܽ?�y?;ew�'�ｯv3�/�P?^㷽C�`��9����>��*����[�����)��(�\�2>U���'0�����=ͨ�>ʎ���X�beI��#>�&꾽g��9���˲�*�7� q��W�쾙���#2���3�H0�:O۱?�g?��&���m��A���~�=I�v>��>�|�>����=����f�]�T�
�>}ޕ>��>���v?� ?$�Ž���?zl�?��>v��j�R��0�=�&O��?�p�,~����о�о�*?���?�5X?��?���>�jݾ�w�=	1�ث?����z��=��*?^�{�\ll?��?�1@j��Ԓ%?�=.>��<��տ?���Uj>�	5?&���z�?�:? �=Z�;?H$4? ��K!��?.�&>�0谽�8ݾ��A�K��9��^ч?����̹�뀿7p)�{�þӊ��K���g�hݩ���	�?C�_�����m�n>�w?@o�@I>U?�u?v��#fy�V����x?�S�WL��t����{-?��w>���?��?�>*���Ů�SY6?��?yA:>'��>�"�=����B?��?:e3?1�>��?��,?):?�D�=;냽ˡ?��v�Sm׾���.z�=ʐw��6�E�ٽ�XI���`�7�Ő�>}w�>~�o�z2E>K�>U�<?Xŕ>hD>H�ξP���v�=��
>�L!>���?i��?�V�?�Z1?L`,?��?�-�?Sp�?vD?4�>��<>yQ?? A�>�b�>�"7��A��K<�I���e�<퐙���M?�0?¸�$�8�qB���>;A?k�پ#���E�1;l>���ߙӾ�%:�������(�}HQ?��{>䀱�DA>��>�B�>�+��ws��E��Ր����0�����e?�u�?~Z?�e
?���>Kt>������?�0�j�>�]�>��^��sV>8�G>o?CMT�����h�{�p�����п�	0��?�j
�>ĉ�=�����K���2>m�?Y.�>�J�>:?�$�<��F�Jk>�4	����?���. ����ܾ�3�>��j?HD�>L��><>�*?W�ռ�����==?a��>�'Z?o�5�b�VL���})��R�>N�s>Z�V���>;�{>+�>;��?�_l?�O6�9�R���1��'?p��?l(��ิ��dn>N�>�6��؇?�:?�T�[���q�k>gT�>Q���S���_�X|>��K�j% ?Y#�>������M�ka8?�����{;��=uv��������Z�>��\���t��Ս��%�=�{:?Y���UD>�>cIE��i\�&��?�����Y?���>��d>�n��[�>LQ���LO����r��>�q������-3x>�Q���ޘ=�"??��>���=����у���=/>����=(�w��1�|?�?�=��E�e��O߇���#?L#��L?F��b"(��X�>�+Ҿ�\�@KZ�'_|��}�*:����?����;�>��z�6<K?/��?Q'x==�	?�Y�= x~�A??�>ӛ�>@���;�o��R�>�$>�I�rM;��/�>�{��0�}��U���r���<�&I]�C�H���u?���>��U?;ژ?z�=.?
�A?�+�?�k�?�(v?u�?eD?���>�?��>��%��>)-Y�,Fl��5��趿���h2Z>fj�>���>XE�>��z?���>��u?��E?܇�>��G?Z >�ƽM�=�-��=$鰾J�.�Žھ�ד��F���@�Ҿk���z����j��{��'J�2:����>���^I�q�A>��>����������MA�}�~���﾿�t�����dP���5���{�>�h1>k��?��>?ڙ?�?:��?4�b��dC?�@p?�B�F �>�{}�$s�=	삾i?,�"�@>�h{��4<��%4��2F>�?�>��>$Y�����?��#?KRZ������̾��w����>�"�<��>���>0�޽��S�Kȓ<���>H��"?&�J�{�B�??:8?���n�G�5
���1>���e =��:�����_P�K�e��pd�6�㾁�ӽ�@�=�n�wb1�41?*:��k����ɱ>�����I�#g�>/��le��j����>��z�~,���Js��r�KХ����=�)��X��:���:>�7�����~�>^��>�ݝ?c�?�&�?���?*�?��!?M��>S
_?[`�?�/�>��待6��ˠ�=,�v��u�?�?P�Ŀ1ڿ`c�>������q�?!-?�w�<�^U?���>)*�?R��>�/���?^�=�q�>�q?$F�>W"�>uL޾����s�������*��>�;7sW>�`���>���!e�YZ���,j�b�??Q�=?��>��������Q?1%>������>�a�/�]?p��>q�?)�>&��>�0�TY��;>2���(lb��KϾ��$��������$��=���
�>mP������Hľ���>v�ľ�")������[��8k">��=Q9;sCr�"�
?�?���?�כ?��Ѿt�M���=�I�>GPk����=b.|��u�"�	��� ?	�<>��D=�B$>��$��K���9|=�߷?��?�p�>On>4݀��>>�p��G>�l�>䕜�D����>AQ>�&?;���>���,c����&?w.�O)���;�m��=�I�?�<���>�wY�<��ȿ þئF??$)>����\>�@վaj0>o�?Ǆ��X�>>:�Q�P�=���=���孼>C�@��!�=;b5�Íྷ�>VP���9��C���=��ھ��?����h�=�¾�߿5����$>�����>T?���>������ƾF�?�"�;ǃ?mᮿ�+v�[�?3�d?`Ͼ:�S��>��׾`|������½-М=��˶L������%�xܻ��\�?�̕=�
d?��ʾ�`j?X3S?Q�?lǖ?�о?ˣ�>7��>��?��>a�^?�?.j�>ﴚ���?)����?Ϭ�>Ȣ�>�6s?��J>��>��/?�1��)x��*e�HҮ�ߴ�?d���l�=�;��9�~?h��>K�8�	�����?��|?��=�
?��?e��?�R?�ݤ?���>UI��n����V�=Vsd?�Վ��PξM4����>����*?'��)=|#>��>.ڳ?�:�> �>�C,?a�2>�-,?di.�s�?}��>}�?N�����>��?L�C�p��H�pD�=���>q����+��C?u�ǽ�5��g'�L����=�Oc��r��Ǩe>�\?�`?iV�>V��>�|Ѿ.԰>���>2�? ��>��Z�{t���H�0��>�=>D��>@G
��9�b�3�קp>��?�=?�a�*`�?�?�)�f=H��=��7��a?wv�=�˾�<�?/E�>=Լ>W�>}_f>���?/l�h���e���8?_��=�N ��E�D�=?���>�v��2.:>�
?��?��	?§t?��>D�>���:�%�ތ:?Dz�=����6���8Q>���=a�`b���>b������Z�;=����Q1D�8��,��棾��
��҄>��˾�f>�i?ɺY��V�\�>iiQ?T��>��D��ʚ����+������տ���>qӾ'TO>&ᮿ��������宾:e9�`"D�OC/?���>�Ͼ��>? �U>�����Z��5?[�0��h���>=F�w>ajf��xe?��9��9 ���>��$?"��>�N�>�XJ�@J'�+>�>�Y�=:�E>BV�>-R�?]�8?�h��,�=m�߽/o���UB�;��<]>�V����@R��͘��O?6Y8?�L
����>��3��r	�P|?��->sw�>]�jM��N ?�Y��M������7V����Ľ-�����D���s�[�S>�t >Ua��Q>y�dV�?\��?�t>���>��?4�8?���?"�@im8?yL ��=������Ͼg阾 ������~��j�C����8>?u���6�=�)�?���>b�E>�GM?w�ξxׇ?.I�>XC?��]?BM6?�Ž�t�=�`�>s=*>���$;�]f"�u7���ݲ��	%>:�<��q?���¾
�y��`e���<j�>e6����۲���h�Pf��k����*k�k8,��(�?��X9�>�����i��j{�?ڦ@`��
J�>a�?r�����?f-�>s��>r�6>LP>��>�G��CD��5v?�3*?�@�?1�&?�h�>�o�:?�I:?��=?��c��5�z���+�4Y��+T�� ��U������?��R?7�?$�D?4|�?��7?6�G���t?ѫ�>^�� �@��?�}9>�rN?�C?�Q�>��v?��:?U�k?��>��?:���I���m.��ƌ>uʍ����>�x�>�td>&��?��=k=�>͋��&R˿]﫿$V�y}i?�-$�,х�c�|���?g?�=b�f�t��>66
�\7׿���>��,��o��Wؐ��ؿ�?�g�����lп�k~?
�=��,����U4?:t?��<�k�=.��?x� <j+��=�?�Vν�v�?����ܾ�/�?܄=���?� X?���<밨>X��;qϰ?�n>SF?��=r=׽%��/(�>�?Lu�?{��=Q	?��ּ��<�p7��%澡p������^/?R�󾘖g?��¿@H���.?��3?&o�rQ�����"��<H���>�>z�ƭ|�������>S��_Z����=� T?�,k?�Y�>�w�?�,?2�>�R�=|݄��)?�/�>o�l?�>?̋��.���O�>�|�|O>�߹>�����v>�|��˺>;F2�Ƨ?`t��5k�EA�XD2?�,���!� ������$)���a>�W?`�����jr�>��>��^�B��<��P<]6 �/��>��$�#_�?N��>��=��>�$�>��>�+r?ʌ�>">�'>�����t�f;�����+0Y����kT���>\}��O7�7�˿/��=a���L,��UF=��=��o?`u�>.h�>�*?>Й?�?�9?���=
�2>�4?�F�?��>$�Q�<��>�a�?�
ȾX�|��>�8�>W��=��t>�;~?�@��#�I�<��ݾ`x�?Yb��s���jN?���?�@n=�s$����>_J۾��s��r�N%,?��?�9?Pҿz��>ǌp?� ?��+�?C&��.?�`Y�p��=�K��`?�j�
=�1��e���v���R��X?h&g�9(��GУ�N�ٿ�Q�V�>��N$��� �וq>[bD���>����0��?�\t���J>�L�?��|��{�>/aN?tˈ>�?n7����>�R�>��F>��g�m d��k���Q?�۲�z�{���>F#�=5���xF���3���-�>9,�ڀ���<�>a����`F?�1c���վ�����#���{?Y'�>�v1=��>gK�q�>@�!�,�-=0�����	?3�C=5��=!�
>)H^�PT��N�>�w?E�9=c D?7��>Q‿Q�>�U~��e��e6==�/=�{?��)z�>5v�����<��>lA�?)퐾#	��[�>�e��2«�������=�ET��˷��d��vN���>�X�<�m�>\��eAf?q�>}ɽ��8?M�?���|�`?]�j>��G�j<ۻMfo>��=F��>�MC����>Ov(>�o>TD���H?#n?��C?�ݔ?T�?@>�?Li�?<0�?N���Ս���f�?�F>��b�d��C:?n��<��>�L�>dս�r�?��J<��=?�������R�"?�dK?"? ]�>s�H=V�D��ݾڡ�=!��'��a������-��������>\qؾPW��G��=)l=try��z�=hĳ?���?�c�=�ic�<g�>��[<��\��Q���>��;>�S��lͼ��_�������褿�A?b|ǽp�p=NS��/n;?��>1�4�(\�D��>���;��f�g<?�&�DN���<�L�ᾰ�?�&��`�����>Tj8?]�?62�(�9���S>c����)�������C�]\�>�.�>�J�����jʋ��4	?FV�C�P=Zq���#F?YW%���e=�wJ�|� ��\ھ}��yT�
�>�J=>X�K=e�L>v�辒X��տ�E�>O��=�k���u���#���>{�>5Y=t�	�o?�E_?g��>�<?$?콉?x�#?��>�-�����Ӿۍ��qy��L�>1�>`6?KIE>����Ǵ�=ٷ�>�9v��L���<�>�8�>?��?��?�2?��w?�
r>C.�n����4�V >�-A?;�#�n-u�;�? �\?�"X�{U��Y�����=�[W���2������@�}�ܽ,:������&�?
Δ>��9?�P��A���C?4�i��9�u} ?�J���2?j��>ɶ�=�獽/�>�Z�>B������;���e>m������=��>���ǃ���7>d_\?��u \>&�>�3{�o��>�޸��b?j
	?"�5�_����>�&?]�I?��_?��?�#�B�
���İ=-.��5�\�徾b�:�%�����C=��-�,O#�_��
��`=���t?���>wN�>PT�>r�!��Z�=��侅����
?2f���}>Zi�<by>�ٗ=#�+�j���
����������"?=`�>��t=���>ٙ�>�(/��J|�c�ҿT�>���=^��Do��x�>��7>�"ּx.׾<$�����I������V>L�����>�M��/�=�{?�'�>6nr�<���T�H�i��Z�2>|�?�>lb�>��Z>�T���;J��w"������>���=���>q<���<?����sξK~!�br����? �H�ý&[b?7�?�|����*��7X�\`��[��3g��E��=˾Y81�P4Q��p�y{�>6G>s6׾�#�>��=��c� �E�޾���?tyͼ�?��Eg?���>P��>�̽���>T�7�̒]=��i��"�>m��>i��e?vmY?�8��< >�UJ����h:<�ɀX�x��?@�<���>[}�> '�?3�'�s����>:�^?v�J�ʯ��jX?�DB?�l?�y�>@�.?��6?Z+��>d�i��b?�ԟ�m�>k=�B,?��>��f�/�Z>#��>Hz�.��<���>\ ���B̾�@�>�K>�4s?�<==� ?es?���?4T���GH>D�>K�\���{˾�ۼ���IY�Fz=T��=/R>vō�k�>6�:y:W��ѷ>k�5�ār?��>�B�ٲ����B��7��Gnk>w���4/��ׁ?!��>��۽�$=�(���} �ؔ��Y��7ٚ��X
?>�.?�9ݻ�rE�6�F?}�.	?4c�?��^`.?4`�>�q��ȉ@��I�>zk���Ž偼�a ��J7?�ru������]��{2i>���!R\�
!���>���=-��B깽���>�=?xҸ>T3�>�9�=U>'��>�
��&����m� >���>\A�A(�j�������I�;��NJ>�>9��>�M.�[���V������uǾ���/ý��9=
�=AF微�g�A%�>G; >�(ս����a�>�"��=��=�-�l>�?�>،?�}�YMK?::���J�����O�c�90Z����f�����>������%��>���"���6���Д�)`<>� ?��F?��1?@�?]�[O��!l">G��>���=
�վ�s���'��y��� �ʿ���Ͱ+���?yK>ߟ\�F�,>S�:?+��9i�>��=��>{�?44>+�������>t|�����e>�����ƕ=��<8�վ�U �1�:�W�|>6�>�����E���D��޾W4�>#��4Y�*?��<��4ҾQً��ES?�Nڽ햂��[�=!D�;m�9?5�2�彥��?�в?��������	��C��o����n4?8 ��HV,>eSL>��Q>�?2�?����o.�mx�>��d>N���>9�>��>�<�>Y*��6��+�<�A�>�y��*�ľY���T>�4��cX�3mV����>o��=���i�{=i�?v\�c�V�\�ͺު�>)�;�8�!�q�Ծ�P>�+�^ه�"���p�4?��0>�G%���Y>,J�8�>��>7;�>q�j>gPɿ�W&?���<��P�p`��o�>�B����8?�s�?C�?�-�>�Z+?�a�?��">���𛽦ȏ=�>?��	����T�7?���>�S��qj�����aC����o�ʨZ>@�>���>E�?��߾�?P13��#��>�;s>���?��P��{�={�r?;��?c��O%�=�ھR�˽sD>�^����ý���L�7>ִ�>%�9�V���V?���>��?=d�>�4/?� I�`�Am�����cU�Y�3�5y�>�	��X?��[>�=��@��E?Ke�?!B?��~��Ǳ���(�6�2��'d?U�M���>84>��J?b.�� ���%��>��>�qP��>�*UL?8�?[f��s�˾���>$�M=������>��c� 4�?݈�>�>Q9�?_��?�E�7w2��뜽��>�*4=���>"/�<���>l��>���>��<@&&>��?���?}�o>)���?r���(�G�h�<�>�޿�]#��v���������?v*���C���N?xN8?n��<���M����F�EC�E县kc�>�l>���>w�R>��?7�?:fV?�D�>.7_?��?�Д>O�8�O�h?�ޡ?=�/?��>F����d��S?*�W��I2�CtG>��>�؋?C+��u�ɚ*?��?��$���B�>� �%�,���L��9�����:�v>_&�>�n>�"����	?v��>3�罁��%�7=�+�=V����?ݽm>sG�=3���A�
�.��ᄫ�Io�����>P>G��?M��N�Ͼ("�>�ǩ>�Z־�Պ>�o<��2 ����=4�������/�b��I=jٟ��(��RԾP��?m��?�CW?K>p?�_�?X������
ܗ���?>Vn�?9��nu˾U� ?�D�?E-[=���Ծ�E�<R�L�&~Y��ŭ ?]�>^����>񫾾�o��F���{=���:����O��>C��?��½[9���]��\u>��>KS:?O�>*\=�o?S�,�s��q��><�z>��e?M�����D��n?Q-�?� �O��~�}z�'S�>9���8�>�>N�F�Fƛ���ٿ&`>�궽v���.��TC�>ڮ�>���<Yx<�7"����\>t�����L? 1��A�=i�<?�^#?��־���6��<5��_ql�b����ԣ=Uо2�R���#?����7�?L���_�+����>P�?�sL�:.��%��������o��=�ۆ�0=߾�i,>����N�?����~⾙1�>k�[?�]���43>�<>;p@��I>Wf�>��>( S>\�?��\8w���=l�?�����$?��t3��R�־&��>�'?R&D?�??JѾ�IF��A@�Y��<xŌ?�#�=�/��?j��?��9�d���3w��v+��_+f�'���$.�*�P><$?߂��?|��>/�Y>�*�>��=GQ?Bo�>d->���>2n�>a?`�>�G��B�Iz�>T��>:}�5���8v.�2ʤ>DD�<�x��n@�k�;VV?
ݢ?s��?��l?�b6?��?�J�R6�>L��4�7��Υ�ThZ��>����I��͠>vm�=�o�Z0C>��[�kk�=�2W>.����w�U9k> �Q?W�>v1�WH�>hg�>O�i������N�e<۾�I���[j�w��+���ti���w=��S�V�=	��>��>��H��l?�݇>3�@=��a����>i!�>�?g<7���u�X�b�.'�����ϥ>ib�C+�j#�9�c�>�=þ�"��@�M�?U9�?j�5?�3�>��ڽ�*8�5I>U4��*X�+�N����Q\>ټ[���l�>&>��!J>�]���5�=Ȯ6�#���
���^�>�l��6X��Ldھ`��>�ھ��'�@bI���y?��=�U1�]�x�� ���I�?'��>�ӿ�)�2>��,>m_?�?Tg7?��?���B3?������?�ds�=��?#�>Zw�a�w�)?�õ��m�>}�w?�!?e�C��ꊿH���0r���	��;V�}K�,���+9��H��fY����>)�Ͼ�O���ᠼa�#>L�<�?3�{?�q&>ܹ&>�|
?�>��6��?��t?-��,�@����;=�;��&>��B�s�9>t�ƾ�3$�}��|���C��/��=�箾��!�˂�!�o�HY�S^��s7?~�޼�*���y�.%�=���>�c�?0�)���?좽?Vߕ?��R?=H1?��y?�,�?����zx>N�<<η�>g`��?����3�q>�]�>sG?bS�>���=&H��QH>��Ͽ����7�dy_=�����Q����h�3��2�&���?��>��оw!?��n?\��<���>N��< ���;s> �����?�	Q>k����о�^=��B�M��>�? 3���v���"B?o-�HY�=�5�="��:A?r��l��>�/�>�j>�����I?�M���Xi�R��5v?��u?��[��(Ͽ{�?��I��c��?��F����?�/��0���k��(�?��D���k���?f����	����=U4r�l��?�ԇ���ݽܯJ�(#�>"��>���T?QD�>7wd��s�?��>k����ࢾ��>�Oս����$�>�! ?�H��^?�ֺ>I<´�<z��?L��?2��?�A�?��2�X:@��̸�?^�_�)ݐ?���=6r�){��B��Uo$��e]��7}��a�)��b�+?��>��?:�?-;P?��ؾ��_?K\���8	��Ǖ�i6)?���kB9>b��'��?�1=�E>��4��E�>w+b>��c>X��Ȩ�?��ڽ�?�B,�ac>a�*>��?�@�����H�����?е���C?���tK��ѿ'��ܴ?��<E�W�g�W�6f�?��?�3?����Ǘ?T:���UC�ȏ���;�IN�?�@W��>�`�=e�ý"��<���[U ?,%+�*�����V?��<��	=�-�a����*\���>�7?��(��f����=��}>���r�Т�4S9?4�N��ƭ��B�<�:g?1I�?���=�v�?��k��
4��?�Ƶ���>���>h�=�y�1)<�E�?"��?nU?R
 ?*p;?������?E$�?+��>?h��cW�+>��=!��I���)ɿ+�>'����?W����i?�-��_��>��	�.��?���l��=�?c������{?���&,�#F��P���6'�*;�><����t�>�͝�o��=�_4�˶>`��=�����V\��X?�?0Y>L[�OIm?�4�?J�>�Ȗ>	�d?���߾��v��W�=��h>/���M4&>搅>��0>4$�>�OM�;�>	�&?~�?�u�gl�=�O�>�f:?�QV�!YQ� �W���>��Ծ����]��?�;C?�;?��8>]�>�ؽ9�y>�E?���?����Ң���C?g���
��>��y�m��= �f>;�[�u3?΃&>ץ��X`F?I�>���=\�F�Q���\a�wi���1���??�o&?��G?���ݾ���>!wE?S��*�;��,��U����>Ư�>�G?�X���8��{�>@>��m>��F?d_��ps�=��?�d�?*�>��\�?���4N%�%Xd>S��<E����s�	qþ�ݾ�b��Tƾ�2��{�ٽ.�|��1�<�Ծ!!ɾ�,���u�����Zr�N��?��O�8?G Q��qS?�w&?9ҝ��i?�1?��L?������?�*>>ݯ�>�BU?i�w?!ᾇXO�έ���Ŀۼ�����a���m���`@��T�ؾ3<��� 𿤢ӿ5����?B|�><��;\S�����>Z 3>�Ί��]�������v��VX���?�!>I?�^���?�;ʾ�ٟ=u�O��g5=�>?�(�R>�w>p��>�k'>:� ?oY�>�{?1��;��9�>�{!=Ec�=��>;����T�>/y2�5}�>��|(4>�p~>l�9@{���+/�>��=�pc�c�¾��
p?��>�n��h���i����?0��=�)�> ��=�2���M<�@A|?k�?�;?��5?ߍ�?(�@�f���=����?�U�������3�5+2�U��?�;A��#�>,��?��+�C'Q�t	l?�%?ŗE��qc?:r:?�v�����̋^��c6��:�U�,����(����}����/?eb羲�ž��?ƋQ?߇=KW@��۵�;(0� �>��?y����o���x�>ق�>�p�=�4�>��Ά4>x��=�8?�Y��56?=e0=���t�<	��4�F?�
@�:�>?C�þ�ܾ8p ����?![o�Q ���d��L��?<6ҽ�+?6��w��?y�K�/��?c"c��
���AZ��5�mQ���`?n/>M�6? �
���R��>������۾�h�2�U> :�>��־<�k?Ƒ'?��~?��M?�t?��a=S_'��Q������6����=ԙ��P־���?�qb�M��?:��� ?�T2?}�;�?Yj�>X�=V��<塾 �? $[��T�?9)�������<>	�Ӿ?�҆F>�
���¾������=(��á�S� �pj?x�>��ྈ������!*@�����A?����@}D�b��?�R=���?f~����׾�b]�*ܨ>jR@��mS��I?ax(?��?�,�>���?j?ځ#?���>��??m�<=KW	?n��>�R�>ۢ�<�ʨ>[~O�s�@�?<߽�r���2?I��J�?r+o�݊r?B��b��?Qq?>9>WM7�.��>IP?I^H��w��[��:oC=������h��"6�_������`AV�@!?���$��x�?�	>�:�=m��=`�E>��e=��߾/;�?�Gb���>��>en`?����jX?d5�� 9��j�?�ܾ�M�H=g>_ᢾE�->_�2�$R�>s$">[n�>1�˾Ǉ�?�]��ܜ5=�V?o��?��+�	�I?�.��3��>8�Ծ��B�Mi�?��j�q�	<�	��{��?�<�ݹ��w<�(T�?�<�Ʉ��#��E�=��� �IX>Y�&���=�i��/ �?b_澬2�?  ���?�*V�������b>xǯ<#�S��KR��D�>?3?_{@;�>�����d�|e-�9UG�ٞ�?������>�?>�%=3��>������lv�>���>��?�:)>b*��΄�$)ʽ��¾��?�?8��>�O?����1�5?7�ݾh+�����~>�r;<!�#�	�>��r?������?KAV��<�?���ԯ?dy��oe=�`����>��
?R"p�G��>���?Žv���n���w�!M�>6�>�J�h^���2?�z?��ɾ�ܮ���U?�P>�Y��Yk?x?z8�>�f��#��?�?	�;l���9��=~���;Ζ��T���n�t�g��Dk���(�Y�?��u�Qq�>��?����F?��.��C���U��XJ>D�>2��EW�>��5>  l>L��>9]�6�>�/��pP
�H�e��l����۾ߚc��h���ݽ$O�?��=�u;>±?7��>Sl�~�����>`Ϭ>��Q>���?�7�X?N�G>�
˾{��;�a>տ�=�{F?�����L������r?7�/?������?�7�>t�sC��|(��>���c���{>����C�=���>�I?f�Z����HEýƒ��m�s>�*���
?��w��� ���徾U�>M��>Uhξp^7��[H���G���f���R���v�l_�?"�����>ى��ez�?�It��m�?:e�����?3@�O�R�iT�L�9>�K>8���~�.>�Gݽ�G�?����X�?��ݿ:7����=��}���?�94>(��?R�>�tƿ�x?z~��5���� ��s�=�{־�A��=����?+�>�&#?|�p�uRk?��?Z9�?��/�\A�v#G�l�=3����q���<>��=�(���B�>X��>d���'?�����'?�8�?p��>c�?Y �>^?�>�C�>�@?�'���
d2��M�=槾P����s+> �@�n�~���ɿ [��@��u����:D���������	��?? �=���2�����$'���f�����%���$B�%I�> .�>21b>��>!�l>=I >��$=�/��:�?�vj���n>�Ҍ>۬�?*��>��ϾTt�<ua����v�V�d���q��I�|+�>��?=k{>V9@?��P?J��?y��&��<�-?	�A#	?p��>��?6�^?y�>��7����z���ݻ"ֿ��C����>��?�>-?����)�?�$y?�ݾS�5����<%��>|��=��ƾ��>$g?,J�>묿��˶>�N?B�?���?�p?GJ{�r_>F��um?*��#ho�I��� @�VQ��Bо��>\w�������P��qTҾb�\?({�>cFv�&�>�[���?��0��Ga�LP��Giξ"+S?��*s��^���*!?��~��z�>���?�H½?2I?�[׿�Ȼ��F�>}8>m9����F����DU)��A?e�?A����r=sh���@?�\��̮�>�5?k�?g��?�'%?+-�>K>5?�8�;�Y�>M6?���;`�>���J�Q=���?L��K�z>˾�S��i?o��>B8R?�U�>��>�ۢ?�?�9?�ݼ��`��3t.?�V�?���=��-?`U�?Ge?�=g?�ާ?�3��$	?�Q���6��M?�S�W5�m�)>U~~>��F?m��?֓ �=�ҿ�>{�6>&�?���=��%��'�=B�;���*���=�콫�Q�55	=Vr
?4H�>���>wD�>�k?�n�ӎ�VN�>����c�<�����羞� ?�2g�G?[��^1���TK��ː?� ��k��(�>%��?:�ξ"�?��>g�0?��>m^p��
?�>?z�Y?T/?>�Q�>���>����˯9�g�J�P�=x�Ub����&��(y?�V���?� h�o=�>�f�=��?��?�
�>ChS�?�e>���>> �>���%t���g�ɂu>���/���9.]�x�"Q��/пf�z��'�9���ƾ>E?��>
�>rR�?܎?Ub�><��>�O�=��9?�>Y]@҆�?��p??M=l?6�>;^��z��q����Cs��rt�-w;��A� �,�� ��>�� �2%?
��?�?�J�B�?�j9��c+��g低(���>��g?K	�%��>�!Ԟ�Y㜿�[��M���.��5�z���m��_\�Ye0���*��W߾BD�>{�G?�7������P��޼?���?���? )�?\Y�e�6��k�*���?־�0�h���k/=?�J=�]>��J���a?	|)>����Ծtn�>in��d�w?ΚV�'۽��D?��8����>SL?6��=T`�h�ʾ�J?�/�w���N�?���a�= L6��D4�x?k���P7?�̾?���d��?�	?��?̣u?w�޾�Q��8��� ?Ip?�9ŽFu̽zk���c����>�x���?���>�����r<?�@?c{;�c�N>y�	��������ϗ�nd����=?~н����t��X�c��?��b?�5?��)?z�?����0�5�@��͌������4?QƮ���?y��> �=�f �ݴ�E(.>Z�?�� ��eȾ>��>d򁿀1Ͼ��E���=zh�>L��=��`?Tv�>l>�`�>�{����?I}?�_ҾZ]?!g@?q�?Cr;���&E�T�>��~�V�/���T16?���>tR�*������(���s�A>aԤ?d��>z�N?X��7~#���$?��s�%4�>F�>>Y;�?�O>	�N�%���-�垈�V�{?am��ar�O��GxF?/{	��}뾿����>ڳ���{���s�%�?���>Ɋq��!�>�>�Q?��޾�>�=��>��>3ʬ�Ng�=-T=�>.of�d���(��?�e`?�7ܽ���>�dϿ�'�>��>�D����e��5|?p�=]�����?��L�6�
��nA>yo�>?)�=�ť=��q�Eܟ?W��?@m?(O�>��=ƪt�hL��H�S�Ǩ��.I���?N�={�*��K�������"�"_�>c�<�|*�?@
6���7?-�y?Q�V��x�=p�1?�H�>��?4&+>-,>c���ð?� �>��>����p5�!W�>R7u>���=+̌��%5?�,P�/�>6�־,K?�Y?!H�?/n�?���?z;��i0`��N� �?�.�V���>�.�?�;��-��?��?M��>�g>E��>	�?�4?M$f�=�?YY𾾪��	�?�ꇿ�A8�.:�����?Bvq�mض=�¾� �>W�>M�M�%�<��?٪�=�CZ?\��?5V\��c�=� �>�S?t'����L�^�;?������?�6��X>��W�`O��9��?�."��e>?�!?89	?�7����?N������>��>�_�>hؾK��PR��i ��m"�Mkx?��2?>5�3����?�'�>~�7?��P����=7b�?��>���>g�:?�	e��]?�W������󎽋F���/$>_�?L�$?/�b=IԬ>ъ)?�C�>�q���˽x:�>"��>�/��s�4��h?�K@��U?�,>��@ؾ��?'?��̿~���k>1��?�x����Y��vo�r�����1� ��>�"�>x����=���>��?D��>��>�o�?�O?{�A�K� �֢=NӔ<� ���[?�N��LU?� -��z�?ȧ�+B����>��`?%V>���5~��U��`�*��;> ��>�n��Aռ�����z�>O�B�Y�$��~��HMB��ھ���=k�Ŀ�s(��<�>�Ys:}^��Y?���>��r?:�9�KV����>�5���1������7<*>k#����*�9��cq?t<��3x��%4��e}?w��o%(��(�>�f�{��>Jh��ϡ>9�>� 9��t��aǾ� �>�L2��Or�kξ�����4?��U?|������^��?�?�iϿ,�r>�BX?�(��X���	���l4��<?��!�ۦ+@�o�>t7�?>���&�,Ǿ�/=GAB�ާھ�X� �>U*�=�h�?����u��������>F��w}_�1�S�<��#���:S�e���새�b�;��p�>߀O�����Ίo�u>%�>�>�k�?b��?l/�ӏw>8}?�Sm?�9�>9�k���?���2'u?�I����e�+��&�<�����>���+���>?�/�Q��&=��+���ó��6�>��>�+?S�Ծ!�<���,>�U���Ӭ=a�9?]����Q�.�?��W�n�>�ҿݯ"?�p?mXs��y�=N���@�y�?f�v?1�E�)o�?ľ!>#@^?�j����@>zZ?�th���>����D��z+j��b-��@�>�t���e�
�L��f�?�>vvx=�[Y��^�=�~
?���>Ȅ`>�sl?LS�r�<>�Fѿ��v���Z�6~��騾M�<g}@>L��s�?��l�����f���>>�ŵ>���=������p?�5?�1_��\|��5�>�t�݁�>։滁"�������� ��Q�C���Ҿ/�ľ�n�?��.?|�K>
��=�z�>rI�>���?��2��Q�ˋ�>����	�>�|�=S%��m6����+�{���gF��{?Zi�=�q�=�Y��z�?�?Uw���>w?ի>����>^J=�w>�̼�m �.����������6â�m~A�����M�?ؑX?�{־)����?�?�ꪾ`���UΨ�ě!�g??1�>iL�?�C�?��?�ܟ?����O4��`��>�	�=��W"8��|d=��>Ku��+�<C%#?��ѽ����BMx�q%?��>�ì�(�㾔��?L.>�9|���!�p"?JB.=鈮>�a�93�?���F>�	V?翑H�������5�).i��O>���>���SU����q?cϤ���U���?�Z�?��%���#����>R�?&�#?փ���E?<��Ψ���w����2�r�*>WU?�m��&o-����?Za&����>�m@=�Α��I�>[��� ��=66�Vl�>Ǘ��J�=�;�>l��?�C-���i?h������=�q���?i�9�Q��>c��S�{�����얼�ʾ��>�~�C]�e����˾��q�a󁾗������$�����=j�����?3�,��t�>�Ӿ�{�?D���)�s�ةI>}�u��1?��?h.�����8+f�jb�= �4��4h�%Ϳu)i��19?�Ԯ<Nx�>!}�01��B���9�>T�t`ǿ��l�����]?=�*?n !>���>v?gY?���>vr?x�?̬��c_���>U�½;得�Q�7Wн64?t���]�>t���V��a�����SԿb6�>y?����H&�>ip|�"�ɾe�����?��.>�����Ud>�Ŀ�!?k�n���ڴ8?�}?Ʃx�k�?I�>�+s�B~��7��?g�?%>?��n��꠿_�	{�/?�篾��?/G	���i���>��ϾB�󿛞�?<+W�'�5��{s?�=��4�?@��J*!����>J h����?J�
��:�>�yy>��>�H���
o?�կ�t�U�Ň8?64�>��?>��? �c?m�t?#\5=邿�@� �>٧�?G[s�왤?�Ȣ?	?$�U=ᬾw޽�'E��H�!����M�kۚ���>�Mk�䋽>����@�Z�3c��B}�>ўW=��k?�Qr��rJ?&�ʿ?Cb���?j,�>��?�q�>��~�(Ľ�����V>�L>x^�>Q�<Ϧ�=��n��Db?�蔾58"�;�ɾً�m�=�W����ƿ�P�?�q�{ԥ�#��?۸��I>�"=�a?�B�>�^P?~�>Sc?9��>`�?J�?�|�>�r�?�ޞ<&�����>��?���?�ս�M�=�u]�R��>;�>?�H���ӿ��?��Ѿ�P@Aܫ?ݻ�?'n���[m?��>L:v?$I¿��(�>: >�p�>T����J����>����7f˿�x������$�>�C��#R��S<��i2����iB4?�?��v>}�!��M?L�7?̹?;�?�ý��������:=(���ٚ�]�b�����疿�F��t�ſ� �F=6��t>;܀�J�j?.�??���?5\?�:��e����?�����=z|Ѿ\&-=�ᐽ�Z>`�>�ŋ>��>h�>������?�ǟ>�mÿ	�ſȼ#�q�$�ɫ�o��>�p�}m?k`n>ʦ�>���k�?)E�?O�?�D
@<��?ν=������>ӟ?M��r�r��u�X��K?jA?�XY*�&�u>���b=�?|��Gǜ>�iݿ��ÿ�/ڿh�B>�~�?o���}=���8��<�T������w����9���ֿ(!H??|{?lh�|��?�������>lmq>�;>�%<?�!?ܯ�>͡����?�� ?�#�u ����?�I��&B� $?�fp��Q$�~��>a!?U�p�z�qf>�$�=rk??�!?r��՘��,W>O`��,2��x>�����>v�V>�5T�l�$<����p>�H_�|ڰ?M\V?FV@����/�>�,��� �=�5A�r�+�N�?��z>��n?���qĿ�罾؆�&g����>?5Sx�d��� 0�� �>��I���T?%����%��l?�vﾫ��:��,9���~>r](>�Z�?o2�?>K>[=� �f��5�>I��>�E�����&>¾�D�JH�q�y�߾�̈́��B����?ܢ�?Sa�=������>�î��G?����W?V>^U�>��N�Q��%ad��}>e�=�¾�8��ڹھ�����辰N¿���j-b��&��$,�|?�!���`0�?G�8��<h��桾�P?cz߿���<����)��3ݿl�d��O? �W�h>�W���?8@�>����M����?h��T�=L�>�:��m�,��Z$��;?W}i�Yv�(��?��ྎ⠽f�;R�R��\��(�?�?�֫>�19���� �;��?N~�>���Un�yg�i��ο�>��= C�B"�ڎ����>�E!��I;��s?�3@p&���Q?�x˻t��Ed?_�/>>@�?1��>�$�؎���T2�@@޾���?[�?Z�=�h�?�t6�V��>. ?�T�=���?Y��>�s�?��?0�>#8V�!a�ė����D��뽽�v8�]ۑ?K�$��̎?�=�D��=��7������2���x���e������n���)�?��f?�!�����>��J�v� ? ���ي>�;��Y�?N��=_A�>���?�V?�Ȥ?�?3?hl?	#�`$i?��H�O�f��o�?Ot�����?rي>�j�> 4'�.[>��>_�j?�A ?��;@�l>�v�>>��=�&�?�@"N�e?�J/��>k����"�.��H���蚿uQg���>@�=|��>�����>9�~?x�>��?�h�>:�=P���~��{�=3d�?V��=�L3?��?�	�а�W�:���?E�?��?���>Y��?c��?:!=?��%?�>�r?��i?i�/?�Ie�,�?oW?�L�?}��P�����>��?&}A��r4��8v����>��.����>�����|�>�|G�4xC���߾�?o�\$$>���?���?⁛��|�Z���Y!�>� �9�g��,�����"8��
?�?3���6;?��v?���?���ȣ<?D+o?��?T�J?a_�
�޾>3�Sv�<v�L���O����1�9?�Zj?1-�~�]��r:?~.�>�=5��='Qx��D?!��>��?j�?�$0���˾y8
?�8$<�H�.�,�	�?Y��>3=�>�e�>�l���{=U��9���G�>��4?����aH��X?�J)��)>�پ}5*?.��>�&ɾP�q?뢚>Eg�>�x�?���{��gq�>hBο�:�?h�Y?G �?�����ޡ?�X�?eп�Z���0�>~��=�s�?m]����
�`���??	��>��?S�=�
�U"��{.?���(��/��b��>\���w� 2?�I\��>F_�?�.�?�0�?���>%.6?d�ڿ\е��1�>��}�˾�?<�>�3��tM���,?`���|�=��?:���vǾX�=�K�O?Z �X�u>������<�&"?F�O>��_?]�<p��i#�E^꾇̤>?�B?:/���|=��F>�І��
�>C����s�As>�Õ�(��s�Q$�?"�ν����B����e��>�%^?Yn>p�R?�X���->`��?fކ=ŷ��f�=DЍ��}K>�c��r�?ʰ^?�u?L��|�>���?'�f�
>>���� >0��W猿�{y�b�Ka���uQ�|���l��>�sL?����`N��?��?��>��>;F"?t��?�F?J��=��*?�~�>Z�;? A��>��ʞ?��>�������f���q�>5J�?ׅ�?�P+?u܂?�:�?�#�?�3�?
�>(�>�t���<��@�=*5�u�
>���?��? ?E��j���?ʼ�>�S��ڄ>j���;L?���>x�?Y?d���>��P����>qE/����>���>��\%>��1��Հ�B�̾��Ͼ�Ƹ<3�N���!?
C���#@�����?G�����=�\?�Ŀ!�5?)nZ>�`�����>����2���iþ$늾U��=/�{�[@�~��X� ��)�F�=��=�_>ݝؽ�w��S�o?_4�]p?��!�=�\���ʿ�|���?�C?)�?v�Y ����?�#��0��B�>�}�1i�?h�=�~D�0�R���]���8?����"пH!u>WR�?`��>j�
?YDӾG�L?Z�1?ʏ����>hz������ھ���?���"*;r�c��ã>��)�.�?�ץ���?OHF�� .?�C?fÏ���=#'�%��T�?5Tl=}>  �?�3t?����M���s�>:N"?�<���s�/T��Ef���-���'?l����Ǿ��>�y'���R�'��>ҕO>���$�\>n9�>�D��d�LQ>��D?��cX�=�)���/��$l��k�?Y�S��>M��K�?��>��L�:8r>�l>^��>b�>�����x��h�O\B��L/�c*�?�#6L�O�����?YF?S�v�
0;?�;?x�ž9J�_�>��f�(�=ڍp?=��j\����߽���>��Ͽ��k���3��T������1?c�>��;??C�NV�;n�C?�	�e���
p�>�>6��>�V'<��پ��˼��$�x��?��>���>�Q?ߙ�?����_x�>8=�?�)��߯��Sۢ?^��?ߨ��L��>Ε?���Q�����>T2>w�?���=N䒽���p����4?,mh?t�?��(?�"E��O��K_�>0i���Z �c��?D-$?2P��pɿG�V�J?���?v�G��q;�[Ҿ�8?Lpۿ��;�N4����=�_?���?�f�?�F�?��=�?,☿� ��@n/���C?��s�Pҍ��"�>_Ha?��7>X�r?B��\�����>ʐ?� �����;O?<�?�+>nid>+2���Ͼ�'�u>�-�?��?O�� 8;�u��L�~�E9��do�莴�zw��߂?~И���?�x��s�>L�e�Α�����t7>N����]?�9��Ʉ���?A�>�5A<�.�>H���4>��P�_�>��־ J���+��ka=KmR���>5{�	��=���?W\>�0�/Q?����?U���1J>�U�>�|=̈́�4d��]�>��5�1ꀾ����UO�/�X�AO:?LQ,=?�ؿj�?!sǽ7�D?H?��?���T?�z(?�ɞ���>NÄ>]�.?�QM?u` ?��>��>?���H��>i;'@������2վ�����S�?g��"���?v��>�s2?�� @���?Ύ���x����>�'�>\��>��=ZW|?q?Kփ<J=�}�澷P�>����Fe�%8!�'(5?�'-?j��<�(�?��0?��I?�=f}^?u�>^�Ҿ�
��@�%?�Yc�/8?Tx�?:��>/�l?#N_?�+?�nb��W��o�>Te?߇��@ſ����� ���m�	?W�>�Y�><[��A��?P/�/ϽFƽі�?k��?Y1�= _�e��?�j�m�|?TA���1>/?,�V<s�e�yG?^�>9������6b?j�>g����M�$�V=1�>��>�>�C�?��@?f�?*v�?�?��?CA*?E>Z��8?,�>Z~�!�������T�2�)&��֨�>����|G,�!�����:��?�)¾�M�%zu�BI?ݑ�>͎c=���/̎?��B�(�e��l�}f�?�n>ݞ��<�ὐ��Z3��,�=�?\�U���>[m=���s�=מg=��v=����4���?Y?O½�b��;ȇ�`t�?���=[-\����?M��?5	��"��?)��?�j�?�\�=�n�s-�>�#F���@����;i�{>��>�-�?'`l?N�n?�ݾ���*��>�Ȳ���>�?w�>?⮙>l�	?�¼<��z?%�>��s�(uW���Z>���>�9�?q&��ο�3m>�>�_�>(�,c��O�w�\�5>L=�qv��W���SZ���A��8���㘽<sC���dᅾ��I?)��?&/`�J���
�?��?mʔ>$h�?��>���T��=7N����>%n�=2�7>դ�>B��M�)�J����|��5�?fӏ��I/?9�>��;5���?X�?V�f��P\?�罐�ؿ���?ڊ�>��B���.�[ͼ�����1���
����G����!>��9�Dȿ��F9پ8	�[�ٽ׭������>T'��w����<�}>�=�>s�>̧?M@@�B˥��.��\�>uƿ>>���;|г?�����ʿ<ɞ���\�kܻ?h�<��P?�=�8�.�>��1���>��j?"���tQ>���%?�>���>�����-i>�8�>��O���2?D�,�l��pZ����z$��pC>dy�>>o��j?�>����>6�&��H?�g#?�Y�����?��?���
�?�7v?ܱ���73�FM? �i��l�W@��Pf���&�w>`����>h/��[�2�����ԾqtZ?�/�>��N��"5?��Y��	f?�J1?�m�M������>)����~�07?��O? ������?S{�>?aZ���=Z��^S���ž��1�"�?yp>�X���:?��P>��?�� ��8���?��6\��QվSx+?��>
��>�r?>�Ž�˦>R�d?��V�l󿦳�>T�+��9ÿ�н'<9>F��>�}ܽ�;��ݾ��6?1�D?&�}��1?J'}>�)J�@�~�΄�?���#�k=��G?ߩ@���I��*�@�1�Z�/?�V��E�8?6�%>V��=�/'?�3��ȋ=&l�����GLk�c��>ǃQ�=�E?������?6���~W����j���?���=|0�Z�>�f?���>�b?�/�=/�N�$����&{�8b�����Y��?Jl�?��
�h��E��=�O�>��>gb�.�l>�s�������ZF��V?"V����e=���jae?��S>�>T�>�.�?�#C?sN0�*�J?�?t�C?�>��>�j�>��=U���'?��?��ʿ�1���Ѩ�x8#>>C1�U=Z>~a�?�#-�g�a?lҐ���%�m+��V�,@���.��c�5��>��>H�{��?&n�>.�>�9���.��[�=y�����?�{>9w�<?�,?L=�?gv�R��>Q�>	�>wY�z����}>\F�<Ҙ=���>��n?|?҉-��|(��
��M�>
�)�4m9�di�>ç���8����<���>�ž�I?b��?�!;?�����b�=Ǔ�eI�>O*��6P.�#7?��?�D��>��h��?���;`��`?A�2?��\?z޳���ѥ�=A��9A�;b�>	T)�N�q>�%��X��$b?փ'��G#>�]=hG���>���?v�?��u>w�?L�?�X?"��ךu>�%*?��F?b����?��M?Bo꿿ڔ��@?�\�?>�>}d;��y?4���F胾۳>��P�{��^UG?���>)��?6T����>2*�����;ﻴ�w�6>D����>���=r�>Y=�l&R��]-@� ��렿L4�?�V?�v��<�:Xy�=/Q>��Z�F�1?�KP?ܱ�>��?K㗿�L�>�^E?r�����ǿBu)?����*R?S4�?��7?�)W>i2�>[}�%'���B�?���>��?a� ���?��?]���B����?S4�=�]z�FK+��QR>�
%��m5�U܉��aC?n?[��w�>q�#g�>������c�0-?J_J?��>U��>���>Gb���P?'�>xS۾��S��ƅ<a��=7���4?j��>s�?;P?�����"?��?�F?�-?;�����>��?JF?	,?%d�?V�#?x������Ӄ�K�>Ӫ�<���ͭV����HJ��ɽ��H����=3xĿsS�?A���;\?���?1����?9Zs?~$ʿ�W�>��о\�����>��J��~��=����S����H�%��!��S���Bg�e���}>x�=!���'V��h?ّ9�wB\��A9�9�ﾐ�-<k���k&�>���Rq����?T̂�iz��f�?=��>��>�5T����>�&9�_��>�uZ?�t?�@>c�3?!ʄ����?���V��?ݷ>� ��V��Y2,?V4���?U�t�`C@>&�O>h�C��D2��?��p*>������z?���1�3>�#Ǿ�a�?>�=<v2=KMi����=��'���"?�D	��
���O_>{7!�ky?�Lt??͓=4n@��q>%8�ӄ?�v�=9ˠ>N>�������>V�> �>���<�혾�(n�*��=}���]�Da�Q� ��{��(ھ#���K�83����н�ܓ>��ԽU69��3�:��"?VvF?��b�d<j��z�>=��>�s�>�I1>�{y>h��������=�C �k0�=�9�����A��þ�#��|�<R=o�eWM����5žO����a��N:�@���\�������욿a����eѾ�H�bk���ƶ��?���A�h>z	�� ����>ұ ?i�;�7?���
 پ�=�F��ɾ�\���Z�vҧ>��=Њ�Λ�{	�>��=.��e���B>�־���<O�u��'�:����B�>�J���=V��>a��>��
?II$?�龳�>1-׾)Ǽ��g���j�r�����?D��z����>`Ȏ>�7��<����>"�-?tJ�����P4X�r���>�=(ϾK��>�v��7�����?Z���N�=��<��=��Ź>D�"?��⾣`i�Z�N>L-�>����c�=<@�uB��",��N~?���>�Cw>�3�>!F?m*?;G*�� ? Q�����4V=����#NB?uh뼨���k�Ծ�è��zn?&��>�r���.>rA�>P�W=�ؾWK�/U��8�?~��>��>��>5�L>�4�=	䢾�0��ٽ�gk>�<?�H?��Խ!����3j��T9�>f�+�Ҕ�<W�3��H�>xGH>�x?���?I/F��Y�7�>��>��>��>�t��=��?�D(�
|">x����ɋ�D���q���=�>�#?���>�O>�?��?u��><L�>���>D��.��&�>��>`'���+>����W�?JF���9�����ߍپ.M�>fAt�2�%?L����5��-<aoV?�3��e��=9��>��M?֘�>ok?o�>��&?8]�>S]����A?1�<cK:�s�>�5m�YoE?!�V�n���+B�<.�=���>;>����j-X>��ݾ�C>�û>�g?M��E�>K�%��Ы�����,��=G����;?P��pk>T�Ҿ��'=��Ͼ��}�7�?���>�o�>�9�f\�>�b�>A��>�*[?�'F?�tl?������z�)�>��%?>^�)?�q�>����^r>�M<?z��>�G۽d'��*�+��Q����{�>�O�>�χ��%>�s��>,������=B���-��>>�Xe�F��>�(�>;��hG
?w����,����>'t���;`>���=<ѯ>k��<m�_>�;���>n>��P�7��>8�����B����=��	>�i�>�LN>r�^>a�?�b�>��?���>"	�?�������y�b�E
����2N�sþ�ᴾ8���C������!� a�>��������>,��=�5j?����q�>��,�9����=��>�v澲A8>D��>���>��F=i��>\�?��=%<S>�@��
�ǽ��?�GD>?��>�yH?��>i��=�'�=gr*?���>\>+�p��>u8���?T�!���׾�\^=J��l^��嘧>����A=�>�Խ�>"{�>���>T�G=�H�`H��n`һ���=}�J��R�S����3�>���'B?wt��N.?��;U���<&������<��a?�G>OR�hU���!>��H>8�>��q>�P#?��(?|��*%N�|�b��0+��P��y��B,r��Ӷ��t}=c��>�i�}&��G;��	j?$��>>�=�X�U�@�]���!?�E����?$�?}m}?��?"�>�#�>��0?%�>S0>>��>�P=�Ӽ>�Ʋ�t�ڽ��`�b�?�o>t3���\�@��=�S7>��>7�s>q�����H�&���ھ%�K��	<�o�۔c�|1C>���O侗?
���ľ�J��cu'���Ήپ;��eĐ����Ra��Y��/>��>���>;Ó>p���멽����=��>`[%��t,>oz�=�'?��p�
UP�����W�>A�#=� %>�w]>%��>IJ��_��>��<�̾��=XJV>Wh�>r�μ��������
?��=6�>c�?U3?To/=�믾���S��;�YB?��>��=1�L��DW>�e���ˣ���h��ܓ���f��ц�
���J+;?��$��t�>۾��k�=Vv���4��O�=�N?�0?ҁ��¾J����S��e�&B:�$�=V�=�+�Ǝ��� �=���=[��>�.�=юl<J�>���键>ә$?ݐ�> a3?>�>y���L�U�ҡ��F���9>s�]����'�=T4���X�<��(��
v��+����㽄A��/`���Vp?x�(>H��_��>ԋ>��p�%F0?�#=_[�Y�]��8?��8?�|;=�c�<�V?�оE�,�r��>@	�w;7��왾�|�>�2�>���?A�@�H�>Z��y���%>H"Ҽ�-�=A^�>��?F_W>%:e=_a����F>ֈ?V��Ƚ�>�)�>3B�?Sq��ѿ��c	�	�޾�|d�y^(��1�b���4�4�&ܽ��>���Snb=:C�>��=�῾|f�=j��-|F��}þHY#>�.>E������<�>g/�>��?���>p[�>�O?{`L?dȨ><�>!�$?҇X>h�[=Ah޾[*i?K�����.>�-���3?��>�J�?)�"8?>�>J�&?=Q$�&:�>&䵾�>ͻ��=
�P>�Z�>������>=?%dc?=r�>rC�>�E?�!=?һg>��d>Hހ>n�>?]��K�~�=��^��؇��H���>0����x�>��羵����@�'�̾竁�rc�>Q{�K��>�V�=���=:]μ��>�~!�Y^�DV龳T�>�=A�d�8?Z�?M?>�">��>�/>��Y>>T?�;�<֒���
��>7'>?�+L>�n�=��{>�l>O�������6Ͻ�A��aGj���~��X�>�H$��?���"��
���/>�oq>�r���>��|><H�>��2>D�D>{�?�o�>�!���?�)�=}�)?�D*���>��>hm?'\�N�4?%=>�	�?,���n->鳕=v�<?OLP��X?��)�M�A?��>��l>p�ɽ��ž�Y�������T�>l�+��A�=��>��>�x?ԧƾ�"�=ʆ�=�X�,0�����7>}=����ˣ�K|��O5j�a��"K$�4��yM��˽k�>	y�aX��g%�>��>4?��0?2�?�M����V���T>bʾul�=�社�Ɇ�����ě>���>�Y�|:�=Y�=۷���G���־c3���>�p���6�=X>2�7=	l
?�z��rN?i�S>-��>1�}���>��=t��>6�s���^���Ӿ���>�F��dW��F?#`�>�YV?��8?�NU��F�>*�_?��T?M��^��>�?��i>�[Ӿ��n��O�<�ۘ�����L�<y�����>������>Q����h?�K�>�t��p�Y�<�G�y�q=�(�= 34��l���{�>Wn�S��?<Rt�b���&'�u7?gVt?�t�=�U��.��gjܽ5�$"���|^>�a5��~�h
>�H�>��>���=̀�>�SM>�ug�)<=r>��k޾a?�s>��7>E> ?�4�=}d����A~n��@L���vK�>C�=���>�E�>��>�Z\?�"=�	��t�gU�<�5нB`��c�>�|e�#�k�^Ҭ�o�Ǿ#�>*��!1<;Y����2�>g!�>e�>Z��x@۾IV>*�޾���^�M�s��;�#���>�:��f��u}�iQ?'�>Z<�?���.2�=���>i�?!�d>�3߾��T��'S>��=4)k������n�>�L�>��1�-'ҽQ���&�=��־�|�q)6����ƶ��&��8�0�#� =b�&�$��N����>9H���`��_��4d\>���۩>�K��׃'����+����5?#�<o_��� {=֧��k�2�3az?^��>\����?*G�;�*��X�!>?w.��&v�`.�>��?<+=�'�A%d��-����>��X&Ⱦ齑=Iž��ƾ�"�=�I��K�_Ϧ>�����D��ѽ/�<��>��z������b>���+�Q>k���>���c���X�>Ef<
�#?���>J��?�K>d����?��>b7�2�
��*�=3��>��@�e\���X�=�W����^*Ϳ��f�����[��#>mLȽ��=��*?�d�>[��?��?p �>�+�=�����YX��s?-3�>�	��#��ㄯ��]>8���hݢ�D�=>W�.?���=�༚�?�DU=�� >�^����=Ms㿲0��a[_����>�?]�k?[8
�K��R?;1?� ?�:?�+��7t�=M�$���Y=)������^>7��N#��LU��;>�)>E�2����#�"�6$�>���=]h>�^�>tc?�@?k�>I8[�,��x)
�g߲>Ԁ?d����I�> �N���>���>:�I�ư�?C���E?��ῥ�>�%�>	i?�%h���8�D0��L��Y�<�h�;?=�>�F�?D�b��Ǟ����?�,��We�?����=A���I? ྰ7�>���>��@��=�?7"�<g}ӾJS��P��=hz��E��Od>��?/�r��8�?`"?% ,>�ą>���?YZ�>t�=>+����_K���=���Jh��{qE?��R?�����A�?f	N���> �������?�@�I!�>�r�>�,ݾ��7>ɗ�=i���f`���?��?��O?��B>�{?��F�Oę=��>vӼ�H?��>BN-�ݡ�>��>�����82?��&���y>��Hއ=,�[�~O}���2�#Z�� �Ꮎ���=��Y?>1�>�l�>���>���>��&h�>o��>b#�W$��d�5?c�?��=x�f�O�>-�)?hI&?��>{�d>ƈ�=�>=�L?�D<?2?r�����w��>��>qs;� ꄾ�tĽp��=�s\?I�߾�S�>*"=��?87d�1b?�\R��(�=�`E��=f?�<�?a��>c�����O>�}�=���=H�;��@>Y��>��o��Ĳ=�z�. i>șU�I
&=���>z�=��>* �?u��>B�?O]&?�������>�ˌ�e��>���>��<���=�pc>�)B?�⣾=ֿA�
�D���j�>w-��:�!��oJ=��>[ʕ�c~ �Æ�?���?z}�����w� ?�9�>uC��ˋ�v{=��>2��>��>�s���1�>��&���w=�����?疃=H5??���4>�	?�h��"X
>k�¾	\�?�����K=�2@�>�,>�L��`����+�8�Z�|?/�>�����^ y�7��Y�z�(���MA?BOB>n������!�G>1� ��w��Om������q�A�����>�ě>��"?��D�Fo?��k?W��a��=d.?�&R��B��||������ޜ/=#��XV�>�A���i$<o:�?�r?�<?
3�>I����)��>�����X��?T9�>�	;���<�楾%��>SM$��Y?�b�>��8>���>�,��5?��&	������k
��Cp����>n<>��e>�%�>���ENͿߥȿ��>y�	>{dz?���?�G�>[��?��?0�?��	�wD��0���Uھ��=?��>5k���~Z�P�f?� �?�)�?�K?u}̾�	>?��߽=�D?oBr��&L����>@A?�v�>�0"����>�%�>H�?%�>ja�>���??���4V?�O'?zO?薏?얀>iKݽkA4�C�=���?3E�?]�7�U����c��\���f�{��?����hΟ>_��uC?Բ�? �Z>��?`��?��?)�=|y>[������)��E?�_�>�&�� �轞�[�i?A���5^�>��?����#��> �����?�����I�(^�>��w��o?򭶾����8�;i�ڽv�+�d�=a�=�E�>{�9��ĭ�:��|��	��>0">�]5��� �Ň�N�վ&t�>�6�Y�?�
'��:�?�M:�uX'?["�<[�U�x�=�î��3���>�v�?W��>\FK?&��|��=���=�N,��Ҿj��>�׭?#N�=aT=�*S�"8�_�z�eɺ�	+����?$?5(�?$&9?�e0���b�������>foq������>�ga�S�@�C?�C�a�e�b}�!Ǽ�5���;��>�7��uh��F?���># k�F����ƾ`w+?���X!?;���8�f�c��>~�?�/>���>�wU���:?f��>8�>�%�+⡽$g~?�\����6��t��_!q>H%���D��>v�5��?�U�<�8(?+���'���$�J�s�>aں�^1 �3�<���d?$n?h��?N��*���P�μh����?�Mپwב�ۃ����Q��?W�B>T䅽��f�e�_�U/H��'�l`˾L����!!>ϱ�? (��r���Q� ���`�#? }�?u�=n����0.��栾 �	>�����4!?�QP����>Pֽ,zp��q�=:�\�H�1?�;�w.?1*H?��\?��}?\l����}�7r=>��?�;?��=n�'�g
�?��?:��>��>^��?��8?#3��O	?�=1?+Y�>�cM>��I6R?U��>�OK����?m�?��3?>�߾�Rm�����־�?�V��@������:�s?Ȋ�g�4?Z�>�������>V�?�?��d>�U��40�>;-�?��?yR��H߆�,>o?��>>2C?�����ֽ;{?X��?�V`=滥�hq�>�{�>�=U�/���?�X�>`Xƿ��Խ�O3��Y���J:���F>�d�iw��s�=�:?V�N?�, ?擬��X	��?
i>��?`��>�GQ?���>��?,k�՗;?�Ľ���=|3�g��?ν ?���>j�u����>�z���?��7��ia��~�>-S?����y)?���=�HM�/6�+8��W۾8�4���>�m�~�>�`�F�#?S&-���ݾ�*>�5�>�=z������~?T4μ(8�`	��?҉�?أ�=G�ÿ,���J�?��.>�G?��������� �>ms�?aHr?eF�'����=�)�>�p~>�x�>��¿Y�<{F?�[?fUf�b*>�$?Ul?���>�9����>z�>����1�Mh�s�0��m#?W��<8����K�?HBT�u>�嚑�1Ț? �4>�H��=k?�\m�s��?�3����l�����;�@�ʾ�_�>���?��^?�h��zȾFĨ���u>��y��Q�?���r��=[L���?f��.=�N��������$�=�e�>�ܾ-�7� ���`�>���>�<.>�Đ>��'����>$�7��U�>]$���D�?�<Ҿ+��?ڈ�>���P������O�?B�?�� ?!g?=���>�?c"�p�#?E���v�o'��
��T>��>�]>�L"��E<3�۽�*?�6�?1!?��]?��ྔ�l��7����`=)>������\���I��	�m�?#�%>U�N>	�?��?�\?���>���>9��>"X?xy�>LOL�3�r?0*n��׆�o/T�+]�o�>!��>�s�=����R��GӇ��#�t�=��q��W��6<ͽȥP?�r��^�V��C�̺R?g^!>��@>Yv�?��7��>R>�
��
�W��?h��>��A���m>$�?�)3�>��n>�Υ>	:�=�B�>���>i�����z?@����޽G����f��;8>-8�>�Qo�;�h�٨�?�?@�`<�T�Cz?P��>����٨b��2U= ��@�>,䢾m-I����O"۽�+4?O�o�H�?Z�*=���>]�⿅@s>,c)>��վ�%�?ׁ��b�A?�d?�!O��U��D@?��?>�׋���5�!�x?W�?�>��
̿\�?���?ل�L����H*<4Ƌ�9k־�p��r�I�������5�x���!�a�5?��������D�G�>|S����Z$?��?r�?��W?f�>�m����W�e=v�!>v�>|F0�� �>��Ѿ�Z�n��T�W���S�����T����n?as�=3�W��r>n��?L웾�꒿���>o{�?�*�?�H?L��==~�?l�L?t�?.,�>K�o�ӾUF?�Y�>�����;Ͼ^?}>|>MDE�bf���⟽`>)�����}�p�y��¿6&��V#9�(�*?��?X��>�Ծ�?=��?�K�?��K�x?3?��+?h��>j�W>���kJ(>��>F�۾Iŝ�m��m���˽ܘ��W����>�a�=��>�?t`�B)ٽ�b��ڸ�<�����$>^j?����?�>� �>��0�¾�L�?|?e�H?���?ym���p[��4_�:��?�ֿU��i�F���¾Ka���#���O�zqľ��C��x�����%\�?%�?���>��?Cg�<�hj��8E>��Z>
A>��M�85P�R� ���.�>@P�=������D�ɿ(�ܽ���f��â��R'����>/4��[�%?S9�Q�n��Cþy2:?���E�>��<?	��>1? K�A��>�4�?��'?d�ڽ�wʾ`�3����>O�ھ!k�=�3?�W��?�JA�)�J�����".P�1@c�ZC?�:>U����Z�>�"�?�K?6P�UR�>���K5�oۼ/�9?�	�??�8?p��D�оt�>��>�X[�:�����!?��}��4���n�v���QӼ����Wm�=u��z^������P��>
>_�a?��;�<�����u�?����������>po���=�n�?�w|?�@�?Y?��>�|�=զ��mA�GK�v��Ϭ��n���>��(��r�>������0��.�׿���?Cq�шc� �����?K?���Ҵ��T�?���>���T.F���?�O�?ˌq?g	b?1O�?�j+��P>������>�#��~��#jc=�K?>�e>����;:�>[���"�>^�?5��?V>�A�><`>��>2󒽝��>wX�>��?�ȉ�N���ܠ��Aྈ���D��y�Ͽ���������>���>�O�>�.�c��<�'J��������?KS�c ��3(?��?�k�?
S���A�4Wi�	����ڷ�wgM��/�=�N>��C�I�k�[�	=-�����[�ϑ��{T1?�b�?���$�i?
�����<���ɿ:�v$?�[?>K����N>e�����G>'gk=����(�y��>X'�Sw`�`%$�+��<cU�>n�@����6�=:�>�x�%��	�>׉�=E=�=��A?c�i?�><͙�m�(��s��(�$��g�2�����R>ږ9��>������>Z�>�)�ܽ/�羻��>b[J>���,�
��Ţ>'꺾)�n����W���b>5wv;%_�>�L?+�Qj���忊5j�g"�yn1>y*?Q�����_?�ey>9w���I�d�>���>�wK?�T>?nl��Y̝���ڿpx��
Z�>q��>�?�BC>��>��=�"�Ǔ޾<�p?�5"?ج�>,T�?f��=�"侹<���6�y!�� �r/����5�c&�>�p��J%׾��\�޵}?/-`?��>�j?������G=���?�>��2��4+>;c�=XLy?nP?�4h>I�3>�ג�(e]���y>fY�>n���E�ľ}������l1���:?69?xJ�>���ܜ>��{���?z߾��D>a�<���z>1�ľ���>��\?-I�?{��?,� ?�'�S���a>���=��>4.^?A� ?z�̿3M��P�.Ŀ�>]I ?h��?��?��x=tC�����#"�����5���h3?D�$?~����͟�0������h�'?���>W��<��=|J,?;�ȼ��>�~�>�=L��|���;�x�!��>�p>���>l2�>b�>f*_�r�?�0�㾶�>�B7�R�3>������>]� ��oA��K�����>�~N>�	U<�Bt>���>X����"]�>cq?��	��T=��?M�~>�3�V,���ٲ?>�P?�N�=��K=���>J�p���>Ls�?P�?9uf�Ɛ���z�^��=�>�9��UF?eYP<�'���C�����.�� ڱ�|�a?�5#<O�(?s��>hS�?޵�?P]B?�)[=n��R���x�>;�� �-?�6�>_d�V���ǿEvN�C���"�b?���>�c<�7o(?�A��_�=]��V�>��>.6�L��>���=���W���]9N�v�=�S��G�>Ok��Kּ�h>b��=]����b���T���?
 �>��῭v½;�����?�-Կ����b����t?p�8>�Z���d����?V�׾AQ3��
?�~?Ԏ-�<�>�b�?���?kwD<F>?��Z>w3�=ն־��켆��=��?W�1��`>���vA��k�>5�>?��	@ح�?��=m9�>��.Z������>�Z,��Vy?,�������y�S�Q��`�'?���?m�?�J���yݽ6|�>/�=�F�ux�>� ?��x>+���ʸ��[�L�(�J�<Fp�;�c>x�n=ř�� �s�-?&�w?��S?V ?���>y!�>�	�?C�>!�>o%��[�W�P�F�ؑ��6�
=NO?�� @��3���0>��=��=�㮿-��.��>F��>��]�RB��'�����=�I�:B�NN= u��'8Ⱦ>�>H��>=��b���|�G?Nw>���=�~���(��N���P���0W=�<�?b�>�5?�lj>8��>TI�?�vt���?��W�N�?�FG?�>�''��A�>��;�@����}`�琁�����$\>�E�>�y1���%?��갾�j�1�?�y?�s8?n��?��>?���?��p?�ɧ��&ɾ=k?��,>-m����>���>)�>��2�p5����'����=O1����?�ј>3�;?�\��xBm?�%>�´?�V�=g5�h�M?5�B?Q��x��>�	�>�(�����7�q��< u�?��>���0���%{%?^�?v����1?�.�a;Z?H.;�������>m0?��?���E��>�Ex��vR�������/�6���:=���>\�>Z���!f<���$��R�=�9���XM<橨>��?�� >��=�灾��6<d�L�Q+��
�>��>5�?z2�=<Bb���ü}����`?u�N?uL�?�}v�$�>\b=K�V�.�Ơ���;a>L�4?��Ⱦ���$��W¾`@;?��m?Cu�?��ܾ��P?w;P��??9�@?6m>'��l�>��?JG�>r�>��=>W��1>V?��I->>�i�L%?Ga>��>X@�;�>fԽF���,�?���9��>Y��>�q?��=52�?�$�?߅���ѣ>w,��$����P^�>;z�>�� ?����E(��9�X������ˋ�iݾ{��`RQ?��?��c� �]?G�)?2#v?������k?�6?���>��(����=�U�$J?Cb�=�=��>�2����T��=_.2>u^��]8>tk ?����Qh>;��?74?i2?�W�?��?���?&��?���?�ϲ>7�X��쀿1�q�>>��;�y�����~�>V㟾>B?ڛ�z8��
p�?ەR?U/"��.>S
���?���h��>Y�>F�D<��w����V��'׼����~X־q��&�=:'��O���?-?('f=;����9?� �=4��>�9׽��վwNf;tD���޻r�N�>�` �>̝�Z� �L,+?���>3����?���=���>Y;����>D�=XO����n?G[�?t�A?�t�>m�'?�Y�> �6�Aڶ���=�_�5ֺ��E����>������?�.*?�	6?�1���~��͟�K�q�?��Ń�Fd�����>�g7��|5>��R�vm�?Uϼ���D���\>��p��Ã?F���h�F?ѐ;�$��?�_�=��¿��7��z��J4��� �>,Q�?�Uy�q� ?��Ӿ�G���;?�sE?Izu=0�?��i?�dA���>�R�?x,�>���>򟄾k�ƾ��,���D�՝h��,�z#��8?���>q����?�Ś??�S�6!?8����>з1?X�9?}nO�%�?��(?�$�=��?"]�>0̟?����������=�"�"0 ?�"?{tv?;铽r�>w�b>�d�75�������~|+��j�>���?UyX�].�n�����o��'@T@���*@�4?מ"?'�7?�T�?�T�����?�>��)�!�����i�B?���fZ��y�d?�h龯�8����>$~�>"�?g�꽻�����$Ѳ�]m�>&j���;[�������>$�� ?��y?Z!U?Ph?���>�j���~��>��Ԅ�������>Nd�?�hӾ�8"�[������>�t���;�����5����`ח�o��lˁ��?�?��?65��E@�>�e�>JKi�Ǌ��קN?G�������m�?�6j?��?s�?Y{\@n?9r���?����"�)��۔`��"?Z�7?`�?d���=����W��⊾�`�>�?�5��s�|�S�P��?��^�͇g����>$[?��@�7?٪S?$iпg늿t$#�������>;?%3}?;s?J�ݾ�Э=�Ϝ���#���e��?ݥ�>6��?�y,����??u�d?�>�x�?���?4I�vn���4�?sE?���?$����4��ǟ�����ջ�U��?yU�?���?�[�?�1U��,�J���f
��nB?eD�>�愼%ǾiR��%�?Y忓Y�?Q�<$�-�Q�=?*�2?��?ƥ��'�r>��ƽ�׼?Go�>�R2�Nƫ��L!?.�Ͽ�e��}6�� �x���j�%�3-�?1�(�����Y�п��'@W%��tL�M��>���?G��>ntg?�i��w�?�3�=��}�?���k9�˥=�R?j�>L�}����5ԧ>�R�>�4�� ��>�ʘ<��2����dp3>�L>������?�n>)NN?``��$0�?R�й��?�)�?�P�T���s�1:����������L��?:���2��ʈ�_���K�?�,P?�[���@���?U�=?v��?U{?䃒?���?�6!?�|�� ��<!�t7?� ��v	��Ǿ�������߿�a���i��J�O?d�?l�t�`l�?���?
����?�^K?��8J�����?�)+�y�
?�iX���p�8�?��ܾ4�п$m�?�V�v����&_���?7	ɽ|`��M@��Q�?J@<>�HO>�q��2�?�M+?$N�?1�?AB�?"���?E��8GԿ�1���Ѿ�f����G��d�=�n?��tX����=Op_>EHX��+���;�>�]���}ĿaZ��~��>_�g��Q��������z?�]�>�u?�ݼ�wU?YNP��?�Ê>�
#>�� @����Y�����+A?�v��v#?�Se���|>�E?d1�$ֈ<�w�&m?�U��V:�?��4>�fɿ��������>���)�#���J?��&?��?��=�2??��.?K�?X�v>!�D;�ŗ?(���m�U��?���?��'�8�C����,�!��?�͵>�?�?J��>:<? ���i��W?�����j����{�h���e�!���}�*?q��̏?df���!ݽ�u
���%>�&O���?�`��P� ����>�@?ފ�.��]��?
��?�sT?���`�?B���`�O?]��?Vv>cM�>�4? �t?	K �?D�>�E�>n�۽�ƿ�pi�	ǿ�檿�<�cی���u����*��>�Ī?o\?����+�տ��&�3�R?�N�<2��=?�?��T?ne>[?��W��OսUV���>��x�M޼�R9�y�.�u>ZW?"~5?�ᅾ�$�>�Z�?6>�?�EF? י>B��>�f�?E?���;���mn>��L�ޠ���S�,p�?�N&?z��?\��>��"�]��?B|�?M�{��>���Ŀ{�?.��O?�Q�kN��r�w�Ҿ�N�?�=���A�=���C�>��@�����?]�?u�?)5���@(��?z�?��G?�-��{^��eq�jEi�=/?�E*��=*<
?&�o����V_�� j����?Kv�?b@#?�|x��<���J���?���>��? n���EQ��i?�H��#%��x�?�
�6��?�ɽr)>���y�>�@I>���>;#?�?I�žߣ��ɼ�ew����O��p?C.Ҿ�?tĲ>̥�>5V�?b��?�
?�=��>M]i���C> ��a�1?n�>�"S������?N<C���Q�!t���B?���=�Ͼ�:��'��>(S�����1�=���^�>H�?C׾������.?�>����?+ "�B�ѿ�Rq����+6P��.^<N�~?��@*�;?~�<%��>L9�����ͥ?g�?���?�`Ͽ��ڿA�뿝�ݿ�&ӿC���>����>�����=�fR?�п�ȉ�ah�>�v�?�N�?��R�-H�D:?s�������f?u�>�M
?w�\�1>�?2k�?��~?���>��=Y�>��Q��j?���?.S˾ T�b���܊?4?Eɍ?Y���Y"�?�!	?j��>Z񣾔��>�%>����Ӭ��GJ?�ž�ڿ��6�\��LS�?ˏ�>��=w*�@U?�a�>��W�$u)?�?��>�T>�i�>�hr>t��!�ֿh
�<�n
�M+0�%?�=DW3�����i>B�ͼ9O�?��u?�k��>̐�u=q?���?͜�?��-?O&�>��1�s)��'9��#�kގ����9���ؿ�̭�=��?/{�?��|?���?�?���>��s?�a��!�U>�?�-�?z3�Q>9>�$�딮�"젿xXȿ�v�=�~�фؿPr߿O�=�=�7���d��Rf?�t=?8I��zr�>�%$?cT��Y��Q�>
�n?Zr��߻���t^?���>���>b:6���>���=qZ�>��Կ8� ?m`?T?�Ԣ�'X�?M���=(��%��=@�?��T?[a�?4Ӧ?������?f~��勿n�ƿ�
�<8�>>a�>n@пd�%��Y��6�q���K<]|�/��>N���?�,¾���&d\�ka���c��Ծ�����8�2�?��o��|��Ќ�J����PпŁ�=�Ҽ=X�@�|=�g?�F�Ƌ;�v�?���D�ܽ��>�����/�iž�w�>�?�����T�>`��?q=��>�c��]���C��� A?��?4���=���?pv.� 4]>���(*����E��?�;5?��T�0?\|1����?�Z���?cC�>�k/���u?JM�?�n{?�ȷ�{�>7<v���F�薿�8�>�/���?JK��Y�W>:꠿	.��0�&�sa�>ZG;!�g?������rr>�?a>�P��r�����E��>l?H!$��6>=�?�!�=�}W�q�D?{�� w���:�&SB��8���ῠ	#?��O��E	��Fʿ��˾�c�o�>��>��7��b��B����z���n?����D�?���?��?@H?�ݽ��Ŀ��=�7�����3?�u�??��>5�Ӿ�T�>y�n���?O�*7���=��?��<�yk>n��z�=`�R�hz�>j�X>&���0ڲ�n3������wx�>��>�CD>�o{?1�@/���
!�?)8N�/��?gN�?/�׿s�@��E�1������Q���?��=�L������3?�1?������xNR?�YW?�u$>�V��y����,?+P�>D��?1&�鄑�v��cz��>?���v�8?�39?(��u�0���?Fו�Vi���Ͽ:Ϳ6�q?6�����.�.�q��BP?]��Z��?����k�.@��:�l�b>�g�?m��>sK�b���0bx?�E>�1�=���zp�o���#�8>�(��4���HJ��!��"6���f?lD?ࣥ>u�?7d?)z�>a�d>a<b?c��>��?N܏?"s1���Ǿ����Ҏ�np�E�=��վJ�r=i�g�*ձ>�j"�k)0?)����:�>���A
�|�d>-�O?�8?d�?w`?<]?9䮽��(�>&�?�vp�cf��f�GC>1S��G?K{>�R��/�-�q����	�;f0*��D��^5�l���]]��RY�.O�[4t�Q-\>H�彥$��K?���>�K�{9'>_��>��?�j���>� )=(/Ľ��+>�QT��p�����c�ŏվ�����]-<�AR�y��=PQu���ɾc>%� �F�>ɂ�</�Y�n�ā�>|�N?T�����w���efR��v�?<�^?=�?}�?Ugr?�e¾f���\Od�E~.>�t��`��Y��R�">w��f<��;�;���o��(��J�]�����BJ>�`?���S&?���??���A�b�b?�k�>}ZJ���9�:�0�ྃ�M��r��| Q?nv��t�Ӿ�h?��b���?���m����\��&�O~þ|��9�&�>�	��i�?��}���>��@��iY��C>�{����?W˽�G�=�9�?�?k��<�j�>I>GO龪��<�d>�E����m;T��Dg��?"'�=����>e�?�e��S��<[ a>��h����=Z�?pA|>�R�<��?ݡ��}�� ?B��?�W�٘@=S�k?V�&�~S��WN���8�o󨿯4]>K"x�-������{���Á>��A��|?)�A�9��?zp>�,�?V?���>��k?jq�>�S*�f�c?';�>�E?�S�>v�?�^L>*wi=���^�>�1>�N��d6]�]�>�����VQ�T��T�\�_�< )�yt�>�����D	�@�@�ǈM?d�p>�?G󒿋�.?��:�>nݾ&��>>62?6*'?q�>�%^>F�+?���6����?��F?]$��gS?v�����>�>N5:�Xf���??&���C��-�>H��=F�S�v�Q��-�>�+�>�����Y?~��?��:>��l�����ǻī��o7>�ʖ>��s�Hq0��<�dǞ��=V�K��?�>>�?��N���ؾV��>B��=��_���V?h%�>�=?�ʾ�w�?� ?��?)��<���?�C���	�٩۾��$#����$ᴽO��>�Q�[�>EC?�:�?n4���?�!о���?`���^?*��w}z?��l�/��).�8P?o)"�i�?�! �3&�>	��`��>:�)>�ֽmľ�k�=م<+�&�̂�����>|]Y��?4�>)J�>�- �b�;?��f�.,m?����X�H>J}�$��>fٴ�l{�>u�b����Et���Pa>U�.?��'?r����:+=7�_��
z;���+���r]�A�?���>�����>�;(?�!ɼ���l�k񥾜!%�>Np��B�=�C־�;�/,�=)y�tsl��j|>˺?��Q?�
?m�>b�w=u��TJ�=�h��Q�fS���ސ��o�M]�>��J>��U?Q��?�?sT?��K?�`�����>��>Ϻ�<n�!=�½>�O �������� ���j���Y�>bQ��(S=J.0?:Y�>��x�#��>��L�)��/"̽�нE��?L	�>��@�Ȓ>��X�~߾�M��H>P�f��-,����>��ξ�'������o>�e�bQ�*Z_=�D5�9�)����Xf���?�/=��a�&�M?�]�=�)*?�]?��+?-׼�� ���;?rd??6�?��>��پ�h��-�'դ��܅�ٹ�>�A?�h�?��H���?��6?SXY�ߵ���K?��#=\0�?�2��⼽��ɾ8�)�Z{�8��>L~Z�ð�=� ���O>��d��O�W��>H�׾\��.T%����>�1��`v���O>���=�<��� �ͼ�=7�S>����{Oǿ�p˾�4>���M�Ŀ���;'s>#G�>��8�@�?=����(�������?@ S��B��O�o�]>i�|��e�>�Pe?��&?{^�?��?�	e?饿>�|�>��>ȁ�>�0�=��>�Y�>��>O�D?ք�=���>��>�O�=�`@�|Z��6Q�W&�m�̾>fB>M5%?1��=���>3��>z��n�?Y�J>��?=Q�:?�?��[��?��'?O����R��n?�9n��kk�>vه>�
�=����N0�����}�T�=��%����?�[@6Ű?�d�?��;��=� ��8r�=�U��}��E������x�o���@���=�w��D�>�.?$`^>�D{�$����Ӑ<5^Ǿo�?���rG>����r܂?#R��p?�$�ޅ�?���Іf�;?_>���?�ޢ�Q9��w��?Js+?�..���=�=?��<��ξ73??=�_?�8�?����!?��>nc�>��.?F6�����?A��Ӊ�T���e�?�(�>�����Ǩ?ܒ�=@X�;����2ݧ�»����>?Zǡ>�fJ>����\]?�� ?�%?�t8=���?���]=\��>��6H��z����>~�>��?���=;&�?ʤ>.��>��>��(?u2L?� )?WL+?ըE?6�R?K�%?I�8?$?i�6�=*2>&�+?Z��=�,ÿ�.������$+?�qѾ��F?ce�>�>�;�ja��O��<ד�=SU��ھ�>�-��`'�${o>�T?�ռ$-!�e&!?'CU>�B��zP��� `3�f� ���Pۼ��?VC���ѽ�>餤�9&t>�p�>��u>�J?ǣ�?�D�>�"?o(�>L��N¹���>r'�S��=�6#>�_*>����Ǳ�E�.v�����=�~?~�N?>!�?�\?>�?_-?�K�>�g�?ISb���/��?�G�?��*�<?�!?a�.�k�%�.d�����j.>�dH�_�H��+�>�w�y`�P?Z���H..?n0���>�('�� ?���dgx�>,%?�빾vq�!r�k_��ϒ>c�>��$�%�>���?K�>�	����>'��?Y��=g_r��P���?0�Q?^}?g*Ǿ�@��{?��� 0>��V���w��H��K,����#h����_&�FkȾv�?�b��F��xwd?dA�>�򨽫U+?���<�?�f3��w�?��>�x$?2�����>�w���q��;Q޾�]�>�%?z�/���a�5i�-��?0?��NS?�m���'�#Dƿ(���jF��s�B@¾�??�h$���?��Q?.�Z���⿝�H?t�2��-ɽ�SY?�7���1��g�=���>��>nf>������?: �L����3�=��6�������>a�J�՝�=V��?\��?o�?�O�?l�?�H�?��=;��?�� �פ�?�?h>v��?h�ɾج@��t���?��������i���P8��Br��\<(�R�h~��l�E�������>�.���>���?3H�>����?�㻮�<n0>���=E荾:��R>>�i�k�`�k�?Ռ���[?Lؾ8��.�?�T�?|��?*8j?��?�S�<�E���>�?�(�>�H?4剾����?�|G��5q�V�������j�j�����F׹�.���RXr=w�������mʖ?��B>y�/?pȝ��f�>C�R?������=�����7q��k	{��7Q=i�����>�g�A���>
n�>2z����>O$�?܂��)�>Ѓ�=~ �>�U�>0g��S���ܾb�&�
~ɽ����>�z?&9L��iѽ'W�>��3?2��*��>Zkm?�>���<J^9>*8?a�%?��B?�!�?S�n<������=���>x�=,y�����ξE\��A��i�ܽ�2�k�K	��!r>��b>e�!�o�M�Z?iz����WzG<�֤?O\�^_��S��?������q>�CD=xM{?��	?�O<�}�>�0�׎��?$ƽ�_��F?������>�����K�(�ҽ�M�>�6���,�&4�=P�?-��=
Ȕ�X��B�j>�_����������=�������`+�>�+?�L�<��>Q�>T�P>�脾E�?�v[���N��e.>F��@�(>FW�>���>�닾�N?���>w���Z>�0?X�>��=%�>Q�s��>�ݾ�o>*�Ƚ��>�lϾ�JJ>���<v�'?"�>��þe~|�*>�>�<�>�t=���2�V>ݦ��v>�[�>W�>���>ʘ�>F��>ž���@>.�=��0>����BP4<�,��H�=�A���>�|�=�>�&�&X�?"��>�<}��r��^�	�6䄽�l%�Ѩ�3������������z�����f_7����= ������>!6�>K�?������ʽ��c>�K����=��J>�_n���>(���}&>
�>v�>�)?L��>/d?t"?��i=k<	�7�,�g�d��>@Z:�0i�>o]�=���;��>w��*x>N��>;�@>x�->(�B��[�.<Y?r*�>�
!?�^�/������<=?��>g�>F�ӽ�Ԓ��\�M%
����?@�[>�.�tٶ>�+����>��C�A�սЛ��a�U��>_���J�>T׽p?�7��`�6�A.?���<�v��X�>4�S>�69��?�:?޺�>����"�#�V�l� ��;�k��J�>ʆ���u)�#Ӿ"����F����<o������ �z:�>ϊ>&C��vþC�ʾ�j��/D��1�5q���оEۿ�V���M���|,R�̀;>^!?��
�@��>���J�"6e��+㾛�>��a>o�i>P-�8t�>��>���>v�>$>�(?�bǾh�>�X>���>O��>5�m���]�aЌ��q��ƫ�=n���	l�=8���#\c>z�%�n���l��Nً��Y��Y�&�q��X���0No>%��>}����I�Ͼs��YB�^퀾ȉ >�䂼�p>V��@Xq=$S="k5< b?�֫=G��=�4'����>��]�`�>@�h�@�>7�����=t�`��#<>�o�����>���=J��������!V���R$�5�?Vf�>&zQ�����F;~>�[>Q	�>��>\�[>�eM��h�=���>v����~�>��n>�>#�̽^T?��?K �>����E���u.H��'��b)���>$~ɾ����Ծ>����(>D�><��=VH,��$����v�웁���-���*窾�c�y J���>[�\=�M$?a�����=&Ե�h�>�"��?h_�2�?�l�!�0>b�J�Ou-?�y̾N8�l&ľ���X�ɽY�<Z1>�Φ=:r���;�~ l����9��=(�ǽ��p�u�����>��>�ɪ�n�?>^�;�%	?k[?V��>�#>��>���'p��4��>�QJ?;�2?s��}���26�A�D���K>vy{>� �>�R=���>�ھ���Ou�>�'��#i~>UȘ�4�/;vP?C��-V$<dMh=�*�>ƛ�>$ai>��=��>)�	=�}�>�}�>/]?�^��*�>&̌>��>�u�<���<s��Ԙ���>&�=�h�U¾N�7���7��0�;��>�����>k>>I��; ��7�� ����� ?�?�5�>e��rD��T�c8�=G/?w���	��� ����E���F��Y��U��p����Wr� ���p�>B>�-.<oJ�>���w���{־�~�A�,?��m�oÐ>�*??���	A?�Q��-��>�m�>�-q>s+
��E>�2������bt>���>�z�<L��><�?�����K�>J���x��u���+k1�4r���A�W��?�о���o l�LR��ׯe�^"�>4��� ���>�����>���=�N�[?W���#>́�>1�6>\?'�;�?�%�=N`?zح�����v4*�tY$��b�=�ʾ�|`��@�=Պ���"���1>� �����0�s'>���=v�c?�u>���>tξu1��ŧ�>m���͑��O>�]������p�=�T���
�1��=��=t�>�+��f��h�gȅ�.���@�=9�>y���ɦ�!>�6�=� s\�e���D=�ꔽ������b��p`<�?YO�=��>w%>w����j�-�y��=BP�>+�þ�/��.�3�=H8?���۸ξ���/c�
�\�0��mѾ��	�NJw�����R;C�7�x�;�����^�O����=�~h��+1��9h>�#�(�=�ؾ��j�~��=�+Ͼy���k�򏾄t[���#�e��>2FL>��	�H.�U�T>������U���><~�1.s>, �Ī�>�h_�i��=�E�WFZ�k�L?7�?�nE�����6TA�����Cľ��!��9?Z�@>}�������#v��O꾄j���Ӥ?��j?�f?����<�c��bYٽ(�Yco��t?�#�ʏڼ�>�q+���(>Byj��X���^�4�L��Ez<��徸�?�(?�"�?�D������vI��Y*=CK澢4B�"U��b�=�D��>�S���?Y�>�X�>3֭�9�d>?%>��>E��=Il??zƽV�?>���;���x'=7�>�Bq���s��\=S+#>���=��>*c �z�4��F�ܪ�<c>c9>@�Z��٫���)?by�>���=�>�?a��>Ceb>�?�q�@=�>fu>��?���ʼ�{0�n��=���"�>L��>��>Q+�#��=��#��)�>���>�¦>F��=}E>@{7>��=9�??�����%��r ���h����>��}=�k���>v��>���毈>%r?^q�&	�>2r>9�ͽb*��	�t+>�y>D\�>U��>1,罻P�i1���>~�>1�Lg��
��'^��MS�=8�`>@�7?:��<ԙݽ\����-?~��>��!�؝�>N�L?Vi����<4vK>�?�L�>�ҽ4s{>�'�?�f��k,X�ԗ�>4\k>��2�������>�Ԑ>��߽�3O=� �>�z���씾oɾ/�>#�>�� ?�T>�P
�H���
�=�)<~� ?B��>��=Q�Z>�}���>�>Fm=�N?���>��>�?=�C�*�!jT>^�>���>;�>�<)��P}>�4!=M�8�C8���>��=��?_^?VS�>�TI>ҽ�>���v�5�U���?��3�>v��J�%>�ʾ6G�>2庽\�4þb�,>�ϱ>�9⾗|>BS�=��!��$��}�>ei>�wF?����
��>M�Y���D?7�}>�K����V=~�(?=6�=��q��]-^��}��>��>�|>��;#�<>0�>2�2?�s��@Bj=]����j?�N�'�n>�4�>��7?�^������nɷ��@O����"?�=b<�%�=r˾�۴:[�Ѿ�g�>Ļ@�5�r�?m�����'�ηB��W^?
}�QH+>��>�P��$??p��T)�>�qξ�C����=�qhO��Zt<���>�&<���=�c����1=�2�>c��>�e0>l�>-1�>���>�>c��Ծހ�HC����>�Z�>�5�>�s?��=�bn�����4a�>�)�r=�a�Q�i�-jľ�GA���^�H����o �t7����3���=e�;>��˽_5���ݾl����oT��:�i�O�9v��]0�=p����=U�7�u�:C�q�U�������s�`Z0� ?�sv�>�0>��5> �e?B���4�w�}��[�U?6�&=
o>7#�={O�oUl���W����>�����ɾk#E��2?��Xb>3�>;ۈ��?�:�-9��	�=@Ȯ=��>&]�!F=��O����>픀=���s���ޒ���n���5=�{>b�z>�o>)�������7��>��>��=�ڈ�
Z�=R�?��>.���	�j�����o"���{>��F{�������rJ�.U?�L��/��?5K>>�d�?t �?��.?����]�5?.S>ݧ>����~O���8��4�4�؂�=�ԇ�)|��},� �?�dܿ	�������>\&ſ�(��̚�dWC?�u�>9'?ӧz=,3?��r>D!G�B��=q�=�e?Q�;�M�f>�]:�L��>�RK;�3�(R�M�?JRa��'�>�oE�\��w���&����3�Ж����?�$?���>=���˚� ����N�?�E.�0(�?x�O?�����%?�[>���>�Mr>R�q>����ɾ��V���>���=����`X�=uo��c�F��|>/?�>ϳ���՞��e���v�>Sҿd�C��s��`}E��1��L��@;=<OV?!C?ȡ�>���>� Ͼg�9�����t�h>�4o<��u���>�:_>�-�=�6���6���?�Ƹ�JvZ�P�U�.�@�g7L?QP�>{��w�
?±	���>��'Y�>4?�~>�:k���g���L�#l|���3�>{x���i�
?���>���>o�>�9N��\�>�c��B�����W��Tž�D�eԾ9��=m��>]��=o����4���e��ξ��(>�ۼ�V4�Ql�>��>;姾6	������}X=�M�/2�>u�8��ž��\��x>>t�!?e?��߾��>��
?wڽA�¾���?��N?2��?+�>p��Etq?�`��j�M���?$,�?�`�=�lɾ'�_?\�>r:���׾<��s�0�7�I��	"����j�D�3s���j;��!>?�V>e�k�E� �;��|=ƣ�>�� ��Ȁ>y�>g���T��>I[?;>��>$�>�V���T �oݾ�[%=�� ?c���4 ���.=:S���Q��;�������Je��ף�=���>MA��Ȝ����	��?[/��S����>�4?m�¿N�>��>�;.?˻>�p��@S?���>����y�F���L?�^>����^�E?8���mK�������>_��}��PF?)�?�>>�j:?�L�>'7�? k>�T??
�A?'�~>M����.I��|�^D��Bn+��b����B>��ᾉ"�wΝ=�Ѽ�o�>,�f:�սwQ�>�"�f�X?3�l?pͷ>ޥ���=���>T,H>�Ϡ?�(#>����Y���I?󼁾� ��yLS�N6*�"�ӿ��G���U�ݾ\���s =y*+���;�?�?}��_Ɋ�S����?T(?v|����ž&! ����~��dH��}�=�?߲��)W���ם���Y>A�J����<��ݾ���>���]��=�<�VR?�X��cH�q��?q)?fo����A�÷P<�#>�� >�,�K�|�l��>r\�1�W�Ѻ,����>�F�>� ��Y��#�<�S����� �L�f"��%���	�rd1>�5	=RH�w_��\>��>
�о'�>]d �Z^�х8��� �����=N��g���ۘ=)fb>��>oDؼ4�e�5�}�Pt�>�I�>��y�(�>�8^�2��q+��PC>������m��>6W�>P@L?�+�?��>ߘ�>�#
?Lx���cT���,�	��ƥV�@�>��p��qx�#����[j�=c��>Z��=���+��>�M>.W=�)>$�>̃�>~�>�\���J�Q�6�<J��+?~G�o���"�qP���o��
�l�D1A�2��Kc=�E#�D�=>h��t4���;�#M��>������8?	QB�����̼{=7@ ���̽Z��>j���]�>8T9?����QI��yQ=4fj?���=�J>�̕�ӆ��Ⱦ��k�#>?�?��P��a�����2W?���:��2����&?�F�=o�>s�g�'���w5B<����>CMȽp����2�2��7�۾��0��M��C�>/���O*�=�[���?a�ƾs�>��?�{v>$ׇ�5�ҽ����ft>�|;�� ���i%����>�޾N����⩾r�%?�{">&��>�?��>=����$?>>3=��H�g
ھ�6��z������#�u>$����?��`-?�2�al>�(������l 4?�2>��>���?[�&��-�vQ�>tS�=d�.�܅��^�_���B�ݯ�Jk�\j�>|1�>�?�>��cy��w~�>1.�?qtϾu/�?�
�?��K�1к>�_u?,]?h��	N>67?���b��>�ӾQ5)�,��D�?�n=��?���>�����6?p�?�|�?��O?/l5?}W"��)#>L�t�$���~�>��=19>]����K�>�)8>}ӥ�I�ڀ�?�O�>h�7=
�G�r/��)O�����>��>.	�=��z�����a?puV����}0c>���>�B�#Q<��=6�e?C�������YȽ5�b?A�=�O�?��?�=�IB��>م�>ʗ�>	�G�^��>�Ɍ>�~;� ��O >��l>���>Ӷt?`2?��}��n�>Z'?e4�?��>˚ �c�5��̶��/�~�m��R���-�>`��o�x���?o�>$��@��+VI?`��П�|W��\��Ca��u�Լ g���O4?pz�?ŀK?�q ?��>��l?)��?W)�>cBN?�"?�ER?Y��>{��?���?G`C?f��>T��Gv�(�W?A?
�i��7�>Gc�?&�%>!C-��1?��?���>*���W54? ��>l2?���ľ`]쾍����+�?=�i�>�NE�x�ý�:ܾТ�:W�y����@sQ�]�����G�Y��ū�>m1�>�'>vㄿ�3D=|���w�>���Xr�?S{?_�@?8痽5|�:��>���T\D�-?9�><����c߾��Z��T=���#��7��V�������Ⱦo`�	�:?>�?�����"?�ג<�=�?%���;)�Y��>�>��r=�E��o�?L�����ҽ�/F�=�>�G1�78k��ѣ��J�����=��g>2š�xc�Cg�?�'��P�����K>s㱾� ��'?t�G?��<���]��!&.��u[���?ME)?F�ؾ�32���w>�@�?<}��P?�E5?=�~=<�o� }a?���?�T���>0
�	lu>3�>64=��>�,��Q>D���+\J��������3˾���fl��é>�u�<�����=ZT���X�~\?<.!?n.�����	?��>͸���@����g>ǆ�<G��/�>�3Ҿ�tJ�cL>�ٖ>�!�?�\�?C����;> .?p��?ſ���־l�
?
?�-v��˳=���Ҭ#��sl���=�2d�$�d�^��>ʵ߾*>�����k��-?A��?�e<?��+?���>�=b4�=2��;6&�Ɓ���=���? 掾�b��0=�%\�=�ٞ?��?�UM?��%�O��>x�?Ys�>TK��oi�?�j�>j��=�ڿ���?5[�=�:�(`�������-U���y����K���A>�?�%��X�>^W?:<L?�}�=aׅ=Pp�>B��>��d?{aj?��7?(�?�=8 ?���>*�0�d�>�^��%C�b��/\W<����d �S��<�=��E?�C�>��/>��>W^���7>�I=5*>3�?�[�YC_=I�d��j`>��>6|a>��־�o�b+��"���ݝ5>��/?%>s?XiJ?���%CH?��>p���֕���?/���fC����˽�{>>6U��ɾGl>[h?��Ҝ�v��>5�@> ��=�ٽ�@�>�Ef?[�ྣ}>���>���;��>�⨽�=`��"Z�~$f�t�~8:���i�=5��>ąZ?�x���U>�]z>`-�?�<�y�A=�#G?����F?W]5�Nb�>Ȭ=�8�<�-;�a!�>6��>��->Q� =�[>�q?�g�>C��{�¿��W=�>�:�>㧯���D�É���Ͳ�Y(N��WE����>��j��r��L��m�?��=x��#�p?z�����=��TY	>"Ծ>mӿXS>�=j>;�ھFU�I��ƨZ>�x�=(�~?ָF?3�q�)?'?�1�?�e�?߶�?X��>7��پ�u����?6O�>�#>��2>"#-�w�z��;��CI�s7�����L�%=K]�@��4J����?�}�3?���\�}^|??�>|�?�7�<��?5�C�f��>¨׽?��>%�?M�)?S��y@H>ˎ׾���>F��>�X;�E�=�s=�����,��������pٶ����������.?Y���p�?���Ǳ)?S�?��c?��w�۾iB0?TN�?��>�Z?	���Z_׾���nS��wZ>� ��R���Ӿ�@վ>�=4C�<,�>|�?6�ͅ-�U�'�{��ȩ����=�?�U���E��:�
�E����=�&�S�?���?J��?j�`?t�3?n�C�eB��F]f����>�&s��h�>N���>��?�L�>�?�6�>��c=��$?pD�>s�i?�;�?yr?T�?"��?S����7�V�~Q�<̊?�!s�xP�Ǝ(?u��<�=fh�>�/?�(���mn��}�?��0?e�$����p~?>� ?��p��C%���?Ȟ> d�?5�?��^�=| >j�?�IԾ-L�>��@&�?�^��|m�=�H�=�{A�v�>b�>
;1����>�V��R,;����D�,¾Vž0\��ړ3>�0�?F�?#�?3�=�c�?]��?j��>�<��k�=���QR?s��?� �����.�?Sc�?��H=]>�j�>+=�>m5?�H�X�]�3s��+�)~+��i
���
����������,�>�s@ia�?�I>?�EN���?�.?��7�{?xx?�E<�e)�r8�?!y?q�?F�C?Z�3?�%���������
?#nD?���`���P?.��>��?�m����>X�S��8?��>w�J=���>�������>눝���
��Q�����?dV�>7�?~T���+�?W�ҽ)I?yM��':?�L?���*f?��?;�(���NZ?�R>�G�?O�Y��NG�&|
?+���)K>&'���	@�ھ��!?�a��=D�?>���?�%?�'�?�����6���k��;��� ��q<�=��$��s���ξ�����邿�p�?�|`�-�>��?1��> x⾇�F�~$�>�`�?u��?�Jo?�?�?�2�=e�*>Z�>���?1�1�>�?sE`?t�4�;;��~Ž�'{���.�'m���>n�}?п�?��?�&j?+k ���?I�?^Ո��0?�_i��T?]#?��5���=�ѹ>�ӻ���2=s�<JG����8��l�>4���;�>~}���ȼ#�̾�|>Kxû���>Gg��?��?f�?�1�?Z�?��9?*(������c>��<?�J=�۾MH�>��>E���9��*����=�M��p	:?6�>?�+@��尿у~=p�:?��>��P�S>v�? ��wD���GR?l-��͚�7�{�����-��RJ��	>,$m?�6�qR�>��&J�uN]���?p�۾��n�v�ɾ������!��"��_v�=r�?�ݭ>�6���/����=�ؽ$_�>���r����`�;m�\>5�<���^�(�h�ܿR�?(k>~\�>�:�?G;>���1V��嗈?z��>_�?��?ʧ?�^���Ԑ?�C�?9�s����?�
���5!>��&��[�ׅt��Q���^տ��V?�F�Q��>/m\�v�+�Y�W3F�4[���i:>tZ�?.R�?�����?ͱ?"�t?W&�>��?�0��у��o���
��>m?/��?J��&�G�:t��?��'?��>\��=��T�#�^�i��俦�ߏ:�
!��M�I>�j�?�$�}�-�����QɿzM���v��ж�$B3�Ľ)��'������wV=Y�Ľ���m���>/���<4��(��� >��ѿa�ɾ�����R�=�1�>�/�Ty�>,??Q�?�W�=h��>�Y�
?�0j���>Dn���?�&0�&n���>`��?[�?��X?���?�1��& �0�@k쁿Ⱞ=���=D�#?�:�>�Q>z��>��A?���Vൾ��>;�����0��\�>�x>?|�?T�?�z�>'?���>CnL=I_�?֣+?3/?s1Ҿ4���4B���9� �����>��$>>��?��?��t�X���3ܾ��?-���6>J���>��4�>A����m>�#n�f3?�|��>�/���ؿ��"�4/��i_=�7%?��|?���>��Z?�9>��$?;�>r��>�b<�`?�!J����ʨ�d�?�D�?Y���i�>�/���ʊ?� ���N�}�3=���>I6X��瀽6U�X��_�?��D�]S~������8?���⃿I*�L��?���m��<<Y�>�|�?��������Ψ<ʂ=��x?��l?x�/\ھ�>&�Q>u$������l>�52�/t�����:Y?�'�?Ij@��=�����;� �b>h��>Ji�?�@?�_����aݿ����S�ؿz�G>i�j?9x�?&�ľ�r��t�?h>�g��U�" ?�Y���/��3��>��#�	?�^D��m\���m")�ĵ�(�����>`�?�ը?��Q=?�);�K[>^��>�-p��.J<�	нfh�Ko@�IwT>�ݽ���?�D��G�}:>Y=?��
�C>�L">��������*F�Î���Bd��N��2���=#,�>�aN?��?��w?�/B?c,�?��D?�h?�?��<?4�A>��>��2=�o�Y�G?��@�ڿ�Fe?�eԾ38>�οt�0��?�bN>�����>~�2�'�Z?�)=.��>�T?�r�2_�����a=�	�*s��t�������ZX��h.���?���>-f�?f�j?�=3?�<�?c�Ͽ.���me���?��޾��$��)��f�pDT���R����a�>���zD?�I�>%e�K$޾<q�=E�-?F\�>7�l���C?_��>�g���>�����@�P���셫�`V��2&?rz1���	@I�ݿi��?�Wo�
�?� ߿Ak쾄:����%�Û���:��`����b��9��	�4�G;��D�]=s��>�ʟ�e�}�_���l�<l,��X�;��?|����t?��>u��1��>K�#=���[����7���
�55?����A?b�I���^�>�{2>��������>>I�e����=U��=��ٽ��>�%�?��7�D�?�D��6gB?h���<.	�J�>�&�����	����>d��ؠ�?���?e������g?Ś �gN��@�="��V��r6?����"�*=�g�>L����ؾ������z���Լ�.��z5?}����TǾD�j�������?�x��k�_>�������N��?���??��;���?�GO?��ѿ� ��3�=�#�>����-�9��)~����(Ҝ��� ���� I<����WH����?߾�>?�}?^��8%,�4'b�$3���P��V�>>u����bq��g���#�>ʞ���h��{BݽAqP?A:��Mߧ��h"��%g����>�8�>��?�5�>]2L?*�B?��n?��%?w5z�����t%�Jk�Y|�>#�9�k�}�Im�;�?�D�>OJ>�؅>
N`?�5�?ՓR?Q�~�0�+����?��?N����i�?*KO�Mo�>�Ո�}��o|�>��?�3�����?�W ����B���p@?���?_��=��I?~挾�{9�S�?�3�.P>�d�>�@�Ȣ���d.�4���]�?j?ҿ�?�W�
�9<+�㿢V�?7�>t>틍���	?��Ϳ�{���U�>x�?ϯ?�pK?,��?������.�?���>�1�>�b�(	?��?����=iC?F��?>�'�}�.���?jV6����>���E/?r���?	?�O>���B��=Z�(@�@?ԟ8?n>?�)m>}&����¿b��?~vd�%*�>�ɚ��?w���eO5@b��>����?�����	M�V-?�Oڽ8]?��?)ە?���=��D?pX�>���=�ǝ>,y&�;.�>!�V�D�8>|sY��}�����1�>?���q'�̱�񍓿�vҾx�0�[��?�<b�Û��=�!�N�?ը�=��?F�M>��>���=%��?<&��ߘ�>_� ?��>��澥
��Կk�\?B���Tӽ,V?�/?י���Z��>U�a��
5?��b�=F�������?s�?�+���>|��?ET�>8�v�?<k0?�-6��xG?˖?{�0>e�>)O�>�a!�7K��E%־1Xy�Y��a��;��=�6
���'>���>d�C?�>�[Ⱦ�i$��0L���s�%��C]�>�Y�>�����靽��׾#�?H��>ov�>'�?�	?��c��0E�&�?Pׇ?�=�t�i�n_0?2-?�C=3�?֊!�y	�� ���{���S0�� Q>y"���=�N�u��Z���|?�+%�W%�X��?վ7�>���>8_?BZQ��b��F#��s�s�l��H��/�@��V�l��>������>�Zƽ`xD=�%�L�>��h@Eu>:�O�P��>���z?��v��{�9|;������>�~�>���? ��?L��>�=����/?/�b�;N5����>x.[��Fξ����2?8�>�?@�,>C@�=Z�潏�S���y�;!l>!4J?�1�?�	�?���~D>��^�)S�>k����~�=��]�չt�iИ>!�|?�� ���(�E,̿�`X������2>/�ƿ@5�;C=�w�>�&3?9�:?��6�E����O(���D�>���?��?U>��K�0vJ���A>xÇ>���mU?6���o����{��#�>�E>l��]�ٿ�/�=�M�;�?->��R��ׂ?�5:>��>� G�)�	�1�0��{?�v����?LT�>A��?ϕܿ<-�>H/�?�>�>��?�" ���c�>�舿Y���i(ܽ�x>��;��R��p�s>~�>?n(�>JAg?���=E��?W�>Ω�(c?�[�?]��=�dT�,�E?���?�����)���s�>���?�Fѿ��]>2GS�g���q5���о�Ba������h�K��?��?F?��	�4پ�y�?
o?D��Cp�?X�9?¨@�J6?ۛ�>��o�3>�iw?�e0?̾��6C>���?��)����K�3�}�n�39ۿAa�?�w�>>�پ!����+@�??��I<2�*?�>>�k��,�\?b�Wq]?r%�?.?龄<?���?�\���?�?5H��l�>p�1�yL>��T�I�X?eѿ/=(���ξ(5>�s��n?�L=#��>EO@>��Q?���?�?��%�y���h֞�l��L9l�-Cɿ�kk��fa����K+��`����>�S?�:���8.>�U8<Gv��㿱��?ٸǽ�/4=�
���6��?Ԡ����H���4?u�� '���� @i�_�-?��V?�|���'��.0��;�>0�0R����>�]?�p�>��^?>�?'$?��1?�(��ܔ?���w�)?f�1�l�1��>_J��~%��k>��>�P�?u�?�ʺ>Yz�=8�ٽ5gi��l��#5>S'�=z�TkW>�=YϷ�{( �·?��<?(�*?oi\?�Q?�	�=]~�>��=Q�;?\e�?�>?[�|����02?��"?VM?�C?8@������U�|�ZE�>O82?��5�|]$��L�zZ>�?�=�w����?v��>�B\��7��4D�>�CO�]ާ=J0?Gb��ۦb>>v?NY ?�s�>�%�>�
v>f_?���>?@��?�@$0�!X!��������*��c�af����>1d-?U��,��>y�>�I=<�B�=�5ż���? @?π���s��+n.>p�����?5��=�xE�r��j���珿����Qӽ�F��R7��D��=�T>Z�:���\���>�r?~��?��>T�f�e��s�>6��v���"�ӈ�>F���?ҿ;���+!)?a�ν��?�@l?g �:�<��H�b�D�-�`r�>�ۯ�K�M����>��ٺ�����3?P�Q>r�m?�Č?~A�>D9��G�?��W?�0�>t�y?�/?���=�͐�;�>���!�9���$���ԡ2�i�<�x�@>�6��=9?��?`N��$����s>��>x�?��t�3�*=���?v��>g��<��?1V�?�Z0�'�?��t?	�<�'N���Ϙ��_�v�>�X�?7�����^��F�I��)�?K��?f�2?)`S?����ſ�Xe�E�̾r�Ǿ�x=�mr��[�=6�`>�F�Q𾾟���
E�>Pm���N�=Sxg��X��=�Y����=�	r?Rؕ��Z���t >�c?�M��ƽ�>�]��Y�?̳�諭� ?�&g?m�I�Ě�*w����?sGD�(�[>�8� �d?K�����>B��><��?����b���`s�l�]�V��G��>�P�c�����?8��>�@�>��)���>�<@�%�?��>������3���S��3nM>\�?��x?O=�7�>��?So�=�)޾]F�?�B?��>�#�z0m����U�=�I׿�ƞ=�x�>ؿ�U|O�F��>�u�?58�>������*?b?ԥ�>��v>@�?��:?��?�ݽ������Ӆ�>��k?׸3��~��ӯ>L?E>�V�_?:�'����?<������&l��ia�?� ��o� �>?ڗ%����>w&?�s1?	a���&?��?�4�>\K���>?�ŭ>R���ɤV�,�?{��E�?+X�>�~���>|2%��ǒ�U�/�ܵ�>�~�?���>Oq��z��č'?}^F�<�M?rOἙ�5��"1��E��t��d��m�>�^���4���`��������?+�?��?f��>^�ڿ��?�D��#\��c������ͦ-��垿x@O#@
f�N����6 �r㶿X�{��W>ۿ��;f���߆�E�K�td��lO�>��w?�pH�9�>��ĽnD��D5��C�@��O�iL���Ǿ����mMN�rG@�� ?�N���R��_�?.�[�/����?0I)@51��0��9�?S��>)h-?��O�39�=6����/�?���>�k�>p昿VT=?j#?�E�?���PR����D@'DK?O�b�(��j$�f���v|>���=�^�:�H=�>rg)������?�%�����?�._��/�M�<p�4=����9��>S�?p>@���>+�^�|���@��7>�a.�9��Ӡ@�%?�\����5��1���?��>�3����?-�?�8�>�o;�M|U?ʠ}�Ig�?xM�?z���;�>��,?�>?S�I�hh¿��3�(���H�B�>��O<S�<�_;�?YcA�w�>vI>EX���	۾L:>�	�>�R_�$e�?��?�G��Q^����?|�f�o0���;��@���>�Y���d����>�����Q�������?q�9?8]�>M܅?d7�>�X�>�?Em���þ<�N?i�i>�� ��{�> �>�����?�"�������^���k=��0=ޕ��v�ؽ�� ?��{?f�?&�|>9�?(�>��|?�!5?!S��,c;?�T��gV˾I��e�>c����b��c���ޡ���?��I� j�UZ	?a3T?�.G>��ɿ���?��s��>|�?H�*��)�>��9?��~=�e�?�}���1�~���"@>Y*�9燾��>�Y�����\�>H���N�<�?*���"���<F{�?>:2?��<�����0J�D�6�e�>�g����=���+?�p�>��z�����?s>�'�= ���]��?���������8?(_�	L?�#�?N*
>�y�>0�D?�?}��������7G:��d?L����ھ/�?�h�?
�?s�ͽee���?����^1��d <Bñ<T�ܿ|����	>�U� ����z��kB�?�����%t��zb�����'?��>�%�>�!���E����L�K�ڽ�B��%�?F����?z���>�\S�O�@���?W��?{?��>p��?�{�>�u&?S#?h�&?R�R�uA@�H)���K�����~�����h=��:3��vп`��r���>�^����>�	������L3�r��?�u4?�9��.2F? Y#?���?)��HS2��V�=|��]?IϿO2�>�?��>k����BE?�3�=�\>;�>�?�����ʳ>��1��VE=��?2����?�ކ�'ݟ�*��?%_���4Ծ��?I*>�jղ?X�w>�Y�>"�ؾ���><5�1u�r�y\�>�A@���	�S3��5���E>�s����G?�e?i濥����j>o+2?Ta$�wD<t�?8ː?׻�>F���������<�E�?�U�?�e>z�N?l��>"g,>ȸ�>�����t#���(�.�ѿ1�?C���7<���?;��*��0��?0����!ѿh$�>�G���G3=nf8��!D�*W;?����e?��L��3
��A����>��_�'��?> ��cʻ���J?5����S4?Zo�?w<�v�>��?�<7��=?����z׶�)��`��?9]	?�?8�ؿ6��?U�j�Ue>��?��>����\��;>�Ѥ?��>�w���~�$?��x��5�����r�F=/��?�8���W¾S5�><���sā���H�����c�?�{ﾯ�t� 2?ְt=�AO>bޫ�W;1?��o?�&��D>>g��.�>ю^=�����>�6f?��>�C��x?Œ�s�E�th ?Lw��f?(;7E���5��@,7j�A�'?T��?;��?F�?��¾�`�(!1?U>X�H��?��:���>miT>�3&=k���p�ƽ����2)��>�<?4,��?k�� ;X�<4�>7�뿭U=���>[7��g�b��"?��.�Ԭ�>�Ⴞ�N;?�~ÿF|��v��>��|?'q���q���F9��#?��>��eT��^=�a���>v>�<���)>X�E��F���o>�Z�<xۼ>�����?�1B?^�j�@� �X��?���?�@?���a��?�>�dC?�ּ�|�rܛ>��V��>D%���?> �?O�R�m���3�u��<������00I?��?Q؛��*h��}>Tv(>%��M�>7#����>�Y@(���P�н	������?�+�>���K?ץ�>F�mϾp���@��8�=�?!3�?��?JŽȧ�?)�Q�"V+?�-�?�ɞ�=k?�
��@>���C��WNx��?T�>ؑ:?ꄿi��.��>�5�>�����M���R߽>�
���$t>W�����K?�O���yq>��w?o�?�f�?�&�>�E? h��P�!�*���i���m���J�ĺ��0~F������:>-(3�6�?��>�>�?r��?�GR�:�>*�V�"=?���t��8 N?�3?�����i��A�?Z˵>��0>�6�>��%������C��亿cԽ=9�>� >`�ο��F?k� ��rE�=�3:?�����/��+?��=�!�9�J��z��n��`�	��B�>n ��]�B�0<5�F�	�T�>տ�>ș-?��?�(Ӿ��v�.�?����6�x����>��?@��>���?�넿'�̾/�?�@?�?�� @i]Կ�~Ѿ�f0���J��3�>R������<��ʾ[�2?�e뿲�??	R�?�y�?����A_��?h>��[>�oN��DU�QYپ��h�²=H���,P9>�ܽ>tM^?E_���?��?ї�?MN�<�?�$���?}��=A]�b�?x�#���3��Tǿ��?h>�>�ߍ?��>l���ǿ;4�GC��)���N�?�7�>+�N?���?�>NS��r+ž�^�?\0	���>gA��z���ڿ���KcC�"�>��;쐔�kG}�vT>�i�qצ=�7�=��!?�Ŀ�4?�z��+_�?Lu���
�?61�>e�>*����Z����(����M��Ͼ���F?��4��3��ƛ��{L�<��N?8k��^�����?�1�=�X���u?-�-�x?��>� ��IP?g�?�NH����Č�>�)7�*�>���1?>
?M�K?䭥?��>�J�=�2>��?��{?�^D��ʩ?�9@�2>EkѾl6�L���q��H3���?�o��ӪB���.��n�>���?m���މ�?bKZ�܆a�'�?
cļ�(�>��ǾD��;R_�u�C?c��?U%?kM�=���=�=��aQ��ǅX=�U����?|_��`I1�\�?oa�>-�X?�h3?1�`��d��y�ξ|@n?Z숿�?E)Z��Bz�?&�O��s���
�<+H>P��>���� )���?���̾�o1?$b迏���W۾��f?�_���L���_?� ?ӗ��ؼ��?=�Q��T�m�>O��?Vb�������h?(0$?�;#Ѱ�_]E>�;��d?�Qs��5=��`���C?�W�^Q�? 1-�ͪ�>���>S���M?�hU�J �?!�N?.ץ�z�
=�Ƴ��:��Cd��/*=��ߧ�Z�O��M�>^֋�B�X?��x?�e? N��@�?8��<�mu=d�ѿ�;?9P���H|�z熿�V���2���>@S%�Yv@?B�н���>{��>/f@�F�>	d->��<K��>N��>2�>�����ᦿ@����!H?��*�>�쿄�u>�?��&=rſ�����?Þ�>8���K���?ϡ����ܾ����$=�-��_U�>m��?d~>�x��DP?a�k?�q)?˯�E��>�T^=Q�|>g
�)��?�=/ģ?����b�����>�h�c�a�r�?�a�=��?!��i�?J˿(���,�g�?�o�8�����4�*�6����T�@�=��A��Pr�}i�[y?ѷh?��? �T?v[?һ�?�X��G�S�8�'���>�g����]�x#�>���o=6�9?M����כ=,\���<���=�:�?�.��ĬѽSQ�>�F)��?�w��P�����?���>��S������D�?qH���L��3��^��?��M��^�?���ۺ>�("@#p6�ŭ�l@��t�?�w�?��
�h)�?ݭ�>�:��i�?[�3���?誾���8?cH4�����?[�þ��
غ������?���>#7�>Q2�>��S?�xq���<��J?aQ˾�J%?�?��|M@>'�w��$�?P��o5�D�1�r�>��?:T��@q?O��>��}�z��>_���)��>�78�F&�?%x
?rcۿ�{��M�e�J���?���$o�>��F?�2��r+K?%:�>/�`��K��b�?�*e:�����H��`(!?C$���W?#�H�[
��	J�����%�?�xa���>ЃB��0ɿ���?�=쿩�5����?R�׾V}<`��?�/?K�?�d����?:��x�k?X�">~�0?\��~�@������+?G'���#�?9>x<u��=l(�kf4���c�S�:l?��$_?�9���>�?{#?7?����o�h?�;�>��?��h�.��v�ɿ��q?v�u?����D�?�@ſ1�5?�������J�C?(7�?�"B?�������?�99�>v�>[�q�&��>T?�^ԾIN�����:�Q�����ž5�z?���{���g�������o?9�6>�J?�N��'V�^o�?��?�*V��Uy�KZ�����o��tF	?�?�>�3;�)��gq�xN�����>�q�w��?��G��!Ҿ�Ȫ?y��?=�=��2+�SM@�,��¤�%�?�u���>��ۿi�t�x���&?ϻ_��>��\j�����7>��>r==���x�?=!��9?��v?~R_=�2h?�Q?W�[?H8?P/4?�F%?Ua?�ĩ����9>��:?%B�>k@;?b>����^���̗�� n?��W������]����?�Q�>�Y5���0��#�?�C}?e���<���!�>3~����z='�������v;�˞�>G6W�H��>�>��ׁ�G-�T�,>�ꢽ��?���G�zd�>#n�>k�>Z6�>I����?��?W��>�|�>���>O��>q�
?�� �q���2{�oa���j�?�N��IJ�>{�u����>)�Qg1>G39�'w��Պ� ?�)�>#ħ=Db�?�o?T�R?�kؾ�ڊ>D�l�Y;n?!�ʽ�T=<��8Ji?�D�><�?5��f"�<"`,��&��$C��^����������@��Rþ$��Cӕ>d�s=Z��2�O>��M?A׾nd#��9�g��?��>xT?"����=�ϼ>��W>ar�$X��k>��=|��UϾ��>��y>.� >�e�=2!�>ش->L����Y?@~{<Y?�W�C��4�}��P">/��<������F?�1?�i?�a?p�P�=1���ɽh&�>��D���X��Ew=k�?�!���>�J��x��>�f��\��΁��[���>�k�>]�2�1>�>Z�	��y����<�>W�&�@D�<��!��c?�F��%��A��=wů>[���ڵ�>�>,[;>U�\���
?��˽8�<?=ڒ�秕��f����">��̽�#�����(�>DY�!c�-vľq��>Q� >WSC>�u'��E�=4A?�3�����O-�b�)?ʥ�>����eJ־�	��f]N�J����j>��J��jͼZ;���?D�u��(�=�����?]K�>��>�ɉ�>����<6����? ��>AV7?����u�>���=�8�>����9B������?��p,����o�U�<�+��i�F�%�	>��>q��>���>Y���JK?�S_�5�@<�7�=��=ذ� �<?)�>t�=���<L($?���������bݕ>
�=׎���r>���>m��>�'����ž<M�>e���E�?��)��ք>1
�??�Kg� ͖��#����"?ѹ��شf�x��G_i?]��>�>>?l	>��>
������=�䌽���>�ԉ��i{>䞽��6>ώ�����j:쾢��>@2;>�n�=�Y\?�O��>y��`p'��&�?{ ?��!����>L1�?^��?_�y��F�D?>�w��Ӏ��˾������e�����'��>������qͻR��?�:���h�����I @ɂ?���>�ؽM2?7;��hH?�@�>Vľ{
�>�>Hk=z������=�A��W�ӿ1���)� > UݽT�?B���W�<�����r�?�\v?:c���?$��?Ä�?�4`��U�>D>��/>8����6�=(6C�(�>�x(�>���r�C�3(�>{�V����=Kq� �>B�a>�=�O>;��>2d�g":>�f���tz>1� �7�+�c=
	�[M.>!���/��>�K�`ԉ��^���C��brG����tr����>�?����Ⱦ��|��>I;����I���=�,�=�;�=c�>>-]�>�T>�q]�	�> ��M��>��y�_~��C,�R@O>X�����JKվUy?М�>Ӑ?��?��E>@���]�>��W��:?�<.�����lK�A�>��,���f����.�>�cs>NO?�8?��>+�̽�+�;���>ӛ]>��E�!���=>Wz=+\ᾜ���yc�=P��>���>(S�>���>G=E���h���"乾M>
�>��ؾܽJ�8䚽�܂>���>Dh½��ھ!����N�ϙ��]!�Z��*�V�*���lF������#��~�>�Mj���h��(�?�"�>u�Q��lX��%ν�?�ا����>[@��-f?K�?�0[>2
���>�?h
�>��]�]�#�C�c��L���#�^�J?G���h�=/%*��F;?I,?��>r������>��>xݶ>�Ⱦ6{�!V��iD޾�,�>l�;�hG�3Cb=}Q=YY��k/�&��g�>��x�7�З��#��>6�>GcL>m'�>)&�>�}�<Y���<���>�3��bm�6R>���n>k�Ͼ�9���#����>}�>'��=r��>4�{j�>���<��>k�_���վ������Ԝ���ǽ�P�TI>m�>GE�<���?�g?�nƾ�� >r ���>�1`���;?z<>-�ri_=(�����=��A>��7��T7�x�k���E�Mx@����>B[Q��=ڇ�<�
q?�����[�>6���!�?&�+?am�>h��>8E�>	dl?:g5?Q�A=?�޾�"�>���P�=?ѳ��'bþ�=��Q;�o��~F��r���w-?&��>c�?u�>?ǾI<���d���M�f�4>��I�װɾҾj��>	�!<�;o���`?t��>3��4�\�pZ��?>�õ����?P��"��>u�ɽZ�]?��^��YD>����%�?s:��,�O������?��Q��i>=��?�޿��2� ��	��?�K'>�:��G�=Xs?�r�>}!��ž�澽
޾�!�-�D>࿽@��=Yp�X��>!L?�c�>��Z>o�??A�?�MY?#������,��&��j�>���}�>�����Ն?�A�5?lQȾ�U�>O�P>L:	?�'���}���<��'��#C��e�>���>Ȓ�>QNR>�V?Vy�>
�?@�\?�=?⋙>��?�&�>?�(?��h?��d?�b?D��9��<�?Q�ps��_ʾ��?1�>e�)�Pl�>�2�?7�?��\�� ���XνF�g����K�6�u��7*�׀b��[�>�^d�5����th����>��=����f��I������/3���k�W�?K�T�>����"�Ti?~���t	_>��G��?_�?���>>H�>��>�HE?&@%?"l\>�)��j�=�X��w?D?�1ؾX�0�v�ٽ�.�>�����ʿ���s�`?i�5?��?�S?7�?+�޾�>o$0�_�?5\�<�;S��V^>?fx>��3?ni�H�>_P��*R��&��;�n����� �6���W>�9>\�>í%�W�>m֗>ƿ�>�Eܽ��<֦�>��?>�ެ�����b��G�/>�,���4�Jz<��V?8��Pb�ɾ �|?�D�>��'��O
�z �>+?QZ�>�.���>���=\�>�s�u��>�X�=A2?���� ��!����^>F���j�J�*��n���߲��6Z?���)�Š���Ú?�!�>�ĉ���=F�E? 9�?K���=��k����Ѿ�ʽQ�T���;?��lҾf ��ѥ?<7?�+n��!2>�H�?��F?��a��u��k�Ӿ��վ���>�?����<7���v�߆o��}?�}f��:���+���=�|>"�>=$�>	��=��W�^y�>�.�=g�>LY&��}�TU��[��>:����B"��}X����jV>#>����]?P�"?ľ?��h��	?�D���u?���>���>��Z�?�A>�%!?G�o�Hb�c�#�ݵ��]d���U���5O�� �>8�>���=#��>f{�>\=���:��>��?��>��T�>ڱ�>��>]�s>�Ծ.��>�rվx�?�e\�;���ŌH���ݽ現���K^þVF>?���>��p?�<?�$?ӓ�>5૽�������=8�x������=��0>�B��:��.k��N>��>�^ۿ"�^�u��<��e�F-��̽m?��w= �D��\��
�>��->� �T`��&�==Au��pn���7�&��>x�e�pd��ҫ��|��>fy�=*�(�.�ƾ��>�u9>==J�Sva�E�f���K�꾪�N��q~>����Qf�d� �K�X?f��;��T`n�B��?;�>��ž��}�n�^?��2?[�/?w��>��>aM�>��? �	>��ھ:�>+D�>H��ttA���?��?{�?�˿�9��1��=�P�<�>��t���>���=�ު������>������LU����?���>ɢ���7Z�_�>e�;�ӹ�PP���lu��?��>����4>�����z\��p����P5�`cx>OV?�~J>Y�>J�?�4E?Ca>�d��*�>譂=pq�>��V=� (�;�����b���ɾ�u��>u��W�뾕>��̿���>�6λ��#����?�Js�3��=oc�0�:>{K�>�u:?��C>�@?�6>��h>�L�?;���E׸�<4�Pm�>����?����~Ѽ�Ǿk��>�}D��S�j.\���T����ޒ��O�����ݾ-y?޹�>�㼸o�=�^�=��>/�㾱r?/�����<d�>�[�>�h�>z��>��:�.��՛-���4>��=&�3����̹�=B{>c��F�R�J�s/�=�!������ؿIꔿ��12��EW���=�>�(-=�C?�wѾ�s>?X�=�eY>���=���� V6����
��>�nͿ�N���#�8>-�X�ԧ��)@��9�>r�(��S��Q��	
]>�,x?z�?��>���>���Ѽ�"k� N��_ ?vq�>Nl?@1�>�>-2����_�����3?��Ծ�*ھN��@?�?�;#?򰣾���<[���j�����fN�@!"��8?f!?t\>��v��Ϫ>_n��$u<�lܼ>VP>>'�>l3�>��-?�h�>��H?��?�n���3~���>j6��X$� [�����u��P��>H"P?�!?�|�=u����B�oo4��?7H>6�B?��;��?��e(*?&x��>2aj�e�w=_'���ھ>�w�jj�<0o�<���?��<�� ���0�m!��_׺%亾H?X6>=O>>�����=�:k�l�?�N�>����y���;i�u2���:�r�>K+?ƝL?'�?>��_>��F��0s��7�>�s
>#��Y��>�n?�r�Ռ9�pϓ�;	N��N��PH���> �ܾ'>HW^�#n{?D�?�,�^�H=��?�>lE?/_��O3�>�)#�KS9����4��>�o1?���<5_	�d��>��3?�҅��P�4n��V�>�6�=����4N�>�n�>���5�B?C��>�?��¾��>��>>��y=z\w�x?| 7�o	�<w����a>ˡT��m�+-<��U���*��Hc���j|��/r��ni�,����n>d� J�>҅d���>�����$�>��PD=w��?�:��]㾦xϾV4�>h[��پ� ��!U���Y��쾌�?��@�=D� ��=U?�b���e���1�=��)?�>E+�?B2��u?Nj?�v��Sh������߾����B��7��A�?�v�>58F�!�,�:���0*>�}�PM�<��2��n����>���>���=N�d>xi��dKX>=�L?g�?���=ӟȾ��.�Xe�>�47�}�U<�?��X1�'�����5��c����E?2��>�2>hb����?p&��9��V��,�>����-f1�F7��I�>V�P��&�?�����	�>g�L>6L?����n�Ͼ�?v�����>�L�>�xɾ��۽Ƽ{��l?�)-?(W�?e�>*�:��U�?�;]�J�P���|�> �>`M�f�ֽ�`+�;]׾= ���?�>�G�?��>/�>��p?a������=ƾ	M�=�7���0������>twھ�"?�����%�>Jھ�b�>�>)�`��U�sL%>�$s>̕���?�A*>H	>�j!��z>�?;-E>�F�=�z>&�g��2��Vg�����׃��c��;���nB��m��u!��[�=6s=��;��p4����>6A�>h�*�;bt���d>�4�����?�h?d$Y>�>�>
��vSt�ڪ��xbz�;<�zKֽ.�O�S���ؾj�S�_7-�§�>�k�?�y�>LF�=��=��+���>O�>�7G?��>��V��퍾��B�}G^����=����ւ�Qfͺ�T=sK�k>B����C�V��=w߾��2���)>lj=4�x�Wxb��	�>��=���>w�|���/!w��T#>�9O�Ư7��"��^|������;�ͽ�>�I�>!�?[�=��r��r�=��V�;�v��|����>�Ga�&��>��?�&�;��>�Y?>��>�*�>s�4"�>�F�=�W@��[?�9�>O0?�A�>Ǎ��e�J����j�=�а�P®��{>ש>�Ҿ>�{n?�=D?���>ve�Z�?[>�Z�?��I?�>zU�>7�?$>`��>DJ�X^=?j�j?���m�~>�?��3��0k��>Gg=�m�=D?3�NM��/��e>��'?�PT?��>P�g�%��=E_5�{K[��<8l������c�Vu�R��=a+l����>�k�����11F�͆Ǿ��/��Ӿ|���"�>n�ľ3
r=Fd���K?�x�>�G+��=��\?֚.=���>zj��h�z>9�߾lZ��q��?�A ��<���?X�?���>��޾^���>�>N�=4�ھȚ�=JQ�=��j��u> І;�IU>���?[M?P�X>��?�u>6��>��J��{�Bl{>"�>���>�U��,���B?Ո�>u��?�ͤ��I>?��>^�?�}L�,��>�˼�o|?{���,>r���)�=�����n�?���>/08?m�5>�Π?]�7?d4y?�m7?:,?��)?�9�?x7?�F<?���>l�2?!;V=	��ɒ>�l?�����廾��>�s?��>����>��!>$��a_=��>�f߾Y����y����9q��ƾ5�<,��f/��h��I轅)i>w�N>�>����K�$>�j�=���=O׳=YpB?���>K(,?���>`�
���#?F�^?�?'�0>g�z?;
�=K��<��?X)ƾ���g�������Y<�ⴿ�{��z���.�gu���n�nry�w��>��W�
~��R�^�#�l�S���޶�d�	?iT>�L����>(��>pkL?�wܾ�)�d[3=�J ?!�'�v�5>C2%��F5��k��:w�>�qI>�*��s����>�x ?�K?�
�<J�>�(�'���\JN=Uxg=X�3>箩=2�>>��߽8W�?�C�>Ũ����TVj?��)�E=p�E�O=Ev�<��>��?�G\\�n���Ph����"?��R�)�r�JD%�1E=j��>��T?�.�!��N�6�]z�v���Y0ľ�4|���>=|�>ϘT����|I?S�p��[־T�?�+�=(��>�G�T�=�b,=G����	 �m6ž �_��`�=Ս<=�$/�M{��(���׏=��h?�a�?�����?�+�=�Y����[��Dl�����>7z�?������d>z������>��@��H*?�Ǯ��!>�1�>}�����>�`��r��A"?���>E�+?�?��+�\������=틈����c��IXY>���s���%�=%/>�_�>��P>_
�>��=4�
@�$;��p?��>-q?ʢ���<j�z�O�?�Ӽ�/�������辬�A��>Ӿs�̼Q��=�@1>�;;>1�Z?K�E?C�>p�Z@�>�R�>���>�%?:�>AU?��Ӿz�=VX�=��޽�V����h>��>�H��¾/��>aF�>??2�>c��>��4>F	o>ĺs>��>�1?K>`?�f�>,��Pgt���}��8��}on=�<���=���<E���;!��N�����z�>�0۽��x?Hg���c?��?k�p>����=��>_'Y?�f;=��?��1k&�͵��W.�>y7$>��=8!�=)�J?��)>Ǔ3?���>>��n�>�e��6�u>ݔ��8z��^z>Ǥ�=���u�������p־�f�Bǂ����*Q�>�p;�����>U¾A��~~�=XN?7x"? ?
4?�D?7��>X}���j�>��H���x����=zϽ<��<����%��>�Xq�:^�����#�����a]�͞龺
�d�j��-�N7n�)��2Ĕ���i��=!;�����
>DQ?�)=%������<
�w=��6=ɴ컂sc����=�RG=�:����aB�=Z�=>/�-9�=-=k>��=���=��=��>�G>���=�0��D>P��=�[>�Gx�<��GnӾD���Y4��C����=lܼ$E�>��r���=_ť��J�>�|3=lz��=�iZ>V��>f�%>�٣>�(m>z�>d�P=�<�gY�k>�=OS{=��>�ǿ�<��9>��+>�0���< v�<sǦ���C�ucC��č�/c������A����� >��!=s�%���<,�Y��*5>�H�,��<��ڽ$��>��=��=�s�=�9>S�̽��!�������=u�w�����Yh��Ȇ�=(��;j3�����qz;��>��= �V<� g�����?��e}$>8��i_�=���q�*>�>��n>��>��>�"�L���������=��a�x�¾��;�n�<��;�Ģ�a��=bߐ��r��	ؾz�J�k%�Iiq>�1�=+BC>[�>�4>p(��ݰ�=��~=���=�y�<,C��k�	=	ӗ=�WA<����=/>�=���>pq��Xy;�Ƶ����<��=2@��']������� >�>>	b<iҒ=��=2�&=���<΋<34��k�=���>,K�=��=��ѽbM�=�	>�7%��	:=�Kȼd�g>/z<f��S!e�7NE��U{��;=�	�=Y>2;��b<�n\<�k>s�ߺ맟�D��;[����~a>r�"J?>�t�;���<bb�Z�.>�����A>�(��y�G��=��7>��g2I�IY�^���y����g�)��w�ȿy��`@��T�< n�<��^����8���=rE6��lѽ���=>��<�^S�^�r>��#>S$=��>4�M>ޮ߽)�L�;����J>SG��+����M>4fn=A!��f���16���=�Rƽ�%�>1K@<2�<�����s>?=�j(�ȇ>��W>CM<��G=x�=�ޏ>7��=�q�=p�0>:݀>]�L�yYN��}߽�>��{�����ٽxC>���<w��%�a=���>���M�>ݯ=X�>=���*�F������>�&���>��B=b��>�Cv�$�>�L�νh�����u3��N���ݔ��ȑ���f>$�:�i�B�=�f^�B[,��ځ�����Ò�r�l>"�j�=�N=�9�� !-�!i�=0q��׍ʾ�o��ǿ>�k��nge�'Ѕ�R+��c���;����z$�S�Ǽ�8�=�����Fe��ӑ�;��=�Z>7G���AA>W��Y�>�St�U;*�����h�����(ս����hm>X�:\w�V� >Y�������*q�2�A=��s<�I[<��^�vg�=�.5>;>�=�'	>��>���k��=��껣]�(t�=��\�(+w>��ɽ�,�;b����r>w��<�� =�.�=��p>�e��yR���� %>[���|62���`�G��=B��=�=���=Vu�=iT_��o�7 ��<٥�;�1���p�f�1��=i0)��ZV�%TW�e�=�Xh>;�K>V�>3Z>C�X��E�<���=��=1��=0�[�~����_>x,���@=>�㽣�=�[�>�i�>���>9�>]��=����b=N94>M�߼���\2�d�3>6�E����2���W ʼ8¹>h�_>�od> ��=��$>Y�g=a��3�6�v'�=�т�;<=���>�9�<��l=�.��м�����1W������-w��1þB�ɾ�嗾R�>5Rx�I�G>�P���d<�諽�9�:�;�$��D.>�ٽ�g���=k� �2���HQ<��u���]>�n�+=F[�<B7>o`�3����0�K������DK�W�:==N�*=6Q��;�Z=ߏ+>rz>$����#=�Ε�׈m>�<�t�YiK�uO����Eh�=�U >s����=e\0>���@=̥�=��B>��	���>g:H���>��=�
E>/�	>%�>9���Jj潔6�<|��<��ʽ�#�A���޶=�O���	��҅=���>��=�R>^�<������=4�<��>��w����=���]�>��>�̎���=f�>��>�q�>ձ�>Ѿ�>U�5�lL�<,"�;�Y ��͵=~L�<�C><K�ɳ�<����fP>:�R����o&���L��qvl�~����=��4��!�/P����<lt(�w#���=x8��[H!=�j@�B��٤��1���X��ҐO���=b^0=�S]�����=��*�PD6==�=���]��-G�D�[; z�>� �>��>�_>w��5=̾[+��#�����>�A*�Ai>�w����=��μ�	Լ`Ѽ��<���>N����W���Z�� =�J�*|>
I]<Gּ4�<��y>�B�����<�5�sr�>&��=��&=>�\�{�>sj��-�=q�>�G�={`����`=��>���=70��>�ka=���>���k� �=��{@��߉B>�z�=3��=��_=d�F=?<=Ԩd>������>z��l�>�F��i���<���}���?�,�>�}l=��>ŃB�D��=(>�F=�f6�m�����W>8�6>�W!�����9"�9]	�O�5����=6Xg�L�>>à�=�G)?��>�>`i>�~$>T�
>���=�uu>�ꤽ���>2H�H�u<�U�f�#>��\> >�i�Xd�=�B�=�UK>u�����>؄$���?�se���x���5��p_�ǳ(��������p���dg=a�>=�ɽ�[���d=���=$�t����;?�<���lW��`M>r<���=๩���i��D�<�U��Wk�/S��aN#>�8S��%A�,;v�=S��mY�'r"���(��0��n�ؽ5��<��Ľ5~��V��<D6?�P�-��/�����̇>%t>O�&>���=�(I>��o=��?<<�B��">�(>��>h����<�7�>�H=4KŽ��� ��$�;�����#2��7P=��"��>��->D>�|R���м�d>���=a8��s�����R<?Ba>�����Uȼ�/3>�e�:�񮾘�ؽ�7<>Mǹ=��Ⱦ�M=t�=!�P>�Jʾce��3�ݽ�.z>T�>�x��̨�=��N�QG<2����m���]=�:��y��Pv�=_y�=�]{<�Hq���=�Tp���D>���=M�j=׊C���<�w<}�>�1@�
F�>�ܻ�(
?ޞ���i���ܽ��ӽ���A�J�;?f��V�}�Ļ�#(K<�ڂ='˅���>�x���_>d��W���������p��X�kԽ��[�b�S��!_�s^Ž0L�=����5V�;7�T��Z�=�ڠ>/Y�>�T>�C>��2�OS�2�<<0G?=��_�!����� =1K�=VK!=)�=�'���R(>�ҥ>*�h>�[�>�U>o��=�)�;E��=ݳ������[�>P��_���o⼡�?�\���@�E�}�N�W�)�־�c���!
���=�d�<ɖ
�j#ڻ�vZ>wQ3>q�{=m��m�=��>�~>A��te=�\�=�u:З��`��s�-���!�wuн=��;�H���.<)J.=��<��{��=�X��>x>)�@>] >0�e>I!�=~�=`��=�.�=K�8;������|�;>��:=��Z�3rD��GY>#�q�i�����p�>�>���ח<a.��s#=w[�=lp�����%��G�>����t�u����r᝾M.�1���@"=u�)������<~>N>�i%<_P�-'<m�>�� =�~�����l�=V]�=t~�������=+��p]T�dS>C%>��=�퐾N�=�^-���>����	������b>��>{Ƅ>e>y�i>oO>]�1���T���c�?>�oW�F,3<�禽�G;>�|����<��S�0|���W���h���;��,�>C½=	b�ǧ���ǻm �����=�߾�>���=��>vܾ���?�?!?FD��ԓ=�ͩ���ž�ڬ��ܙ��� ��b?�N!�g�����ƾ�zۿZvR��ོ����g�>�X=D>(?9�?�����R�V?�̮>���?�5m>[싿�>�����9<�Vv?�/V��Rt<�|?�h�+�?��Y�еg?]J���Q~��i��e��>���?f��?꾦>�6>v��=��<?N욻-67�ѕ���/���>?p@r�4�Ľ�_]��)?Y�ξ���>>ؾ&�>?�D��A(�2�����7.�Տ�Z�$>L�V���-?
Ⱥ�d�>63ھ�D�?4�P?S�?��ξ!d��q?`/�>T�%>XA?���<�H���O�JJ��[�e>X߾8�=m��"�Z?L�!>{�ž��>sA��XZ���k�K�/��������>������x��U��d ��se @���?	.G?h?3c$?d���M=P�?��0�w�ľ��v�9�=8eW��!�V��9�?�=C����h>��%ѿ0<8>Q]N?_��=~ 8>�y=���=ɹ
?L�ݽ-k�x]p�(p�>Ӊz��ؾb!п�d=�f�ҿ%�@]?��?�Y�>�))?|����>	o��zs���T���B*?�����/����.���Y��S�U>2:�p�U�iSk=�]��U?�P:>�m�>�g>��4�w߭?��=	b��'Z7?��->� J=4��w"�"_e�F�,�C``����Q�>_�%?Nr?6,?�Ɍ?��<�M?�?�\ɾ�Y?�.���>?��?ُ5��
?*V>9� ?+�#�V�>I�?b��?g��=̿�#,�Y6�x���ú;�kH�>C���A��gd�ڿ�=4~=���Ƚd�M�yo!����=�L��'�> �l>(7�?K m��
T>�?�>}���F��?��/?���>� A���H>�ؠ��]�>��I��K0k�d��a��=-/?1�L������?&���'V/��<<��<?��W��Hm>�v�3�?�󈾢��� N����?�?s�i>�ԅ>�qE?�|?��� �u�^�<��g>jM�"��Ad��5�)�?I퀿]c>�b��Ε�����"�?<S>��H>֝޽����Oh�[�?٣�>��?j�t��V>�D2��^羪?¾7���>���cS�G�Ǿۻ��j?YK���4?IYs���?�K�>p2?E4X?���wv�>��r?�}�>V�>��?81�=�þ>&�����=���>�g��+Ⱦv�U��ƿi������>�Vþ������>k'n?���,?帕>�E��������>0,,?	e?_?��ǟ�=/2
���^��Η=��Ѿ#¾2C�>���=��Ƚ�!���d?Jgr�צ鼱�ſ�>��>׽S?��{���>[h!?�x�=��??��?(�1�?��ٺ��ʕ��b�=G
/>��r���=?�Xy�_�<h㊿�	Y������q6>��>�$�>M�>�:�=��7���
?N�#���4��z�����>�.:�H�{���O>T�#?�Tj�~��>R�Y�͚
?��W�1ߙ=��>R��Ӄ9�:@ʽ� �������?\w@?�=L?�׃?ɇ> ���k����!?��X=��p�,rw�� >H}>��9�XA�bu�����?�W�?e��>��d>��|=��>w�>b�>�E>G�?��#�i�����_�`wL�u䅿�� �2?�?_ %>C!?Z�P>�	?���=�*�B�{?��>�6;� ?��>��,;b�>�O�=��ݽ:=�����|�{S�>���m�I�>�>}�=���>��~�H�r>!�����>q�i��5�=��?�'��Oۈ?򲢽���=�)��� �>�T�>}z�>p����>���>p%b�ah{?�i@u��?���LM̿V�Y����4
��@>��4>˖����_�>?�{����=��p? =��@}<;?���#,{��G2�ܵ��I6`?Z��>v��UY�<Vڀ>���9-����O�Q��>�3�?�ž%�D��e?M���\�L��ػQ�r?h?��>'�Ծ�$�=di4>�q׾Ji��;� >VW�9z>��`��G4?;ü>Q�>@=�=��.����Z���'!?�B�	�g>�&��4?�Ш>V���Ʉ�8�?VP�?�(?30�>��>a�1>�Ⱦ� U?�.$??�>w"�=��M=>V>H�Z>& �>`/@;��?n߿DL �p�]�S�J��/���ɜ=��	?G�=�5�G`g�X�?!$ɽ�k?r�=�ʥ����>��:>;��>z#9@��?��V��I>�Qq?��½0�����J��>�ǻ�dQ��N�)>Fܵ��z���-�?��?��:?�խ>^3;3{)=Ze�K`��>��>��&?P	{>�}������G�!�7�� �?}�a�� �?�ܾ�n?���b9?�Ԟ?^��?�;���6��ZM?+�A>���Q!��_?��*�J�{����Ĵ�?Ax��*��Y��)u?;�=.31���>�����f�Z�?h����@�o��Hӈ�
��y� �0�������=�ў>/W?ք���:Ӿ7g$?y^n��-�>�@���?�ݛ��������p�!��> n�?�W�=�E�}{%>Ĺ��xF��{!g�U�#=7R�?4��?�y��M�|�ﾾy�>kb�	=��'?�v>��>X(4?uE�?�0�?�Tx?�?>2!?��?��?ґC?��>vԑ?P��>ݳ��i&$��f?�?�.=��M��b?�r��\��;>H+$?�4?5�y�N@Ӿ��M�jH�>!�	�XM�=�J]>�����=ǆ�>�I8?YG&�[:�;�tT>-Ǔ?���>����i?V�>/aA>\%ھ��ǿ"�����־�j�=\��`�?�n{=6��? ��xx�; E?Ͷ���f=��?m��>C��>�"W>��>���9���t�bp�-����|��+?��׾�����w�dr�?���?��t>A�?g�9?�z�>(���]뫿�� >��!�a݋?zY��_�?n�Gb?6So�v� �_�v��`0=��l�=��Xg��X��9�žu��=��!>�@~?�h0?O��>����<5?δ�<?$6=x�g���>]u�=~ν��h�ӆ���r}?�I^�ԚP�/�?ȱ�?
��Q��>:	&=,{G?XmV��v�<��>�l�?.|�?�JQ����<��>R�����q?�#{�
^�=7��9�V=��:����p_���R�u�/��j��� �
�>>9'Q�e�?������>�?��^� �r*!?�7����?3ػ�����9T�����@�ԾM҆�Fp���Z�?!�꾪�	��˱>�4/>��V�܊p?���>��%@�������P�����1��>��>�_I�6�p��C�>�t=w�X>�x�&/�=���>�!l����?�>�~�<
��>؝����>�u>w�W�
�G��䩿��>fw�>�܆��B�>&����5';>" (?��t<KO�>�=ξ��/>�;�?l4�>	D5�=<q?<�=��O[?M5N�Ս?�?�N�?�� ��O>O�}��N��������ʽ��[g�,sB������>G}�>���>�,�>$��>��^?y�ּ���>/M�>��{�lh�=�����I۽������㌿�:���^P?�=�����y��[&�������@�<@X�*?��>@��>8,�>�'j�@�q��;�?]e>OW?�ɽ��>��.��>���ޏF������{+��8I>_0���5���Nl�_?*�ھ�j�>]�Z>�`?f�z?ϳ�>[�v>�ݙ�������JH>��I���.gB��a���
���=��>Q�R>��I?ג>�e<?�F�>�?_�?Q�>�;>{� �Wo�V�����&���`�����qI?8�3?Ґ��<?�1�=�i>Z&�=vc���?��P> �?r*?+���M?�2�?ySw?��������;?i��s�8�+��%0�'>�����|_>&vW���s=�99��+¿$�T�򈾬	�t&�80?uY���� 0¿O�?�*���<���L�׎�?Tk��#?���?+U?>�ߎ>���m	��M����D���ϽL-�>,e=3	?�� �S��?���?Hp\?���>�V��7�����@��"�>+�7?m#��8Б�H�ҿ�վ��L��J���a8���� �!��
��B���CV�_�����>�2m>�"����v>�y��+�=�5?�O�,��>���=q���?�?��7>d�7R�>�e�>9A'�kD�����>�I�?U>�?������c�z�><���(��/���uyy��X�?�F>im���籼K�V?0�پ�u�?���E@99�d0�c�>^-�>�غ<E��=���>��?$Hy����̴���꡾J' >����G��9X>>��>IX������?��������&�|���!?x�<>��>��?W�������O?�>v&H>�[�?��?oM�?��P?3�������Z���=��3�����C5��'-����=�[���>�������[�F��˾
��>8���r�G?y��>.�1��{��tU�0Bÿ����J�>��?����ݩ?�p�>�����Ɓ����?�b�eT����>�L�;�#0?V�W?��i=$	���R�4em��+����> �>/.�?�����i�>?��Ӹ�>�/N�*j�>�����>ȑe?Z�D?'Q�>��U=6�X>�퍿 �?T�f���i��y{�x�m���5����>�
<=4�?6��>-�=:\H��c��D>=}��-�>���?��&>R��w
�>�,�>��B�2f�����=x=�g����V5>i'd=���?��*?���{�8>���>�@��m�
�]+���"�>����\�.,?2�?7+g����x��?�.�j+E=Uj?v�5�\5۾�qɾY�>N-?��|�la5?+N�=���>1�&�����>SY{?Ţ��k�o?e}#>�J��s�徠ǯ�v���ݾ@�澙\�?[6�>�M���,<�?�Y;~3���c?�)�?� ���>{����bw?Ge�>L�R?�8��̄?%է?��¿X(�ZVC����>�H����ƍ>a��>��u�U"��XUB�ʌ�=L�?�E��?��G��F�*:>A��>��3��>ӽ�T���H�2X���O>�d���M���x��)ִ�@ꕾ%�����L���?��̽�|�>��澦�P?Ƴ�<��-?�U��m3>IA�>&;�>8�9>:_�?GF?���\�>f_�?[�7>"m�>Vn?d�*�lJ��޿��V?�ҩ>��<�羯ѯ=x<n?��
�i|.��T¾��>(/ؾ��F?w!��D>��=�|�%��:9��?N�X?�N�>�z�=lё=�{$���?���NJU����S�\>@#,�����̚�B��<v2��$_��Ax���C�>��=?�8q?l�?�9?�M����+���,?S޽>�I�=�ѿ��i��i'?�/9>��e�X��5/��k?j�Z��:3���1�<�>�|-��%��x�>P]�v���SL���.=�^{��*
?D�Z���H?���.?L�>Ne=�Q`���t������jF?/
.�$�>L�?�噾�٫=�c�>a���Ȫ�>סF�N�`�/j�?T@���=�x�<��Y>s�|����>�G���ˉ?X3�� �o�������Q?=�T?����5�^������>W�����7��K?�@�Ⱦ����ܘ=�慾n=?k�>՗�>�ߊ�l8?� �?�H�,�v?�^����I>�SY>�f>�\��%����t��:�=�Bc>;�:>e�`�/�=@���ގK���&?������>�����쀽R�־�LC>f�?OB�>��N����?�i?��#��H�?��>�?]�q>P�Z��˾"��>U�����?�*(?��p>�G���s�dR䂿x ���Ġ��S?�3�=bú>��>0�%>��:�����V6?dǅ>[�׾�Mo?P3H���>P:C?.���;�/�_8����n���=��p�	ꬿ� ��@?�y��Y;��&�0>��m>_@&��n9>�ƈ>�'I�=0�>">�Y4�޻>Sz:�O}��P��w�
�v�����^�r疾��?P�O���+?h�*։?6%���Mm��ة��	��.��?Hj�����ܕ?��>��|<>�!2��,���>k�$?f�?V��>�3q?kDE�&��>���j��=��j?J?��G�E��FD�eD]� �"�3g����ؿ�gc?��t?^���	C�%�?M`�?��K�����)39?�n:��x�}^�>���=-�G���@)�X��%=�͎Ŀ5�?�2��R�n2?�Ԍ?GΩ��(��@�<�Ȑ��k�?��d?�&f?W^s?j\����z1�>�����˴�S��>�c��ξ:/���c?�S8��{"��<�� /}?BW�>�_,���>��R�pb����?(�'���?��&��?Ssݾ�������?K�?;����>=3��)��? R�=��(�Ⓐ?
�@� 
�����u?	��m����j*>��2?����-;�$�0�V�g?R�>羢l9?	Q���̻?��g��Ͼ
�=LR��?\B�?��>42�?���Z+O���Q� 3��
B�?%\�?n5�?P�g�n�R?W�?�d��L?E;q?��N���?<S�!v/>����ܾ���>���>�B�>��>?o_?��?��?3N~?3�9?ڷk?;�g?�&?��u�rp?�/�>��?�}�>�h���A��?NJ�� �L����]�?.Ys��Ȅ���I/�?���YDο���>>Z?I��s��j�C�������=7�G?�,?8����c>�(?���>S��� 0��b=��$>^0"�MF�>� ���H�?��?�$>��h��� �gz�>=�>��>�?�qR?�PC��8�\dX��"�?�7�|���%ތ�}����??�P^>�?�政�5@��K�=
����>?e�Y>_b?�T�?{��*_�A?��ؽg��=ew{�@�Ծy��^V�>]r>eI�?���/Z��a���%7�=����?8?��5���9��?�@ן�}�'��?���5�޾����O?�
d�N�M?,����Y�����3@?�I�?BҾ��>=��?V�[?����lτ��b?,�t?~n���+?�pt>�p����?*ͻ\5���=���=3E���)a��Ϛ��v�>|�t�9�H�,��:w�>*rA���m?+U�D禾,"j�&=�?���?t� >ZC�>�H^=V���>{@�
'?�^�?X�����
���>v=��	�ߤ%?�7:��? ξ��>��??�t=F {>�̃=�D�=�ǲ?�t��+��Ϡ����>���>N~p>9�=�J\r�~$�=:��>~/"?�R���?ؾ0>���>����Kw?W��>�0?�G�<��e?�;����e���?��a��?��{<~���?��=}&���t?l
?�/��QW����>�y����>?�#�$w�?�{�?��H�^XI?#/?g%ǽ�_n�>�M?Jx�?��>�o�Of��lt��� ��&ݾ\⏾�J_?�9��}?b�?V�>�LU?�>o�?��Q=|�A��A?8���H�=M��?�OY�O�z?6���k��<���[���_ƾ�[�����f$�>D�/���_��&�>����m맽�K*?"DK>��q�����zC�>�i?��>}�*?�M��\�;�z=N
��I�3?�	?�Do�g�|�6Ga�պr����?����?��>\D�k�N=�?-�S�$�=��罬ʺl���S)���q=����[&������M�=���>���>\�C?5�ྑ^�>l�"?$�?G]�e�?���>.�=�5O�"���E?"�ʿ���=o�D�M&�Β`?Z� >�`�?��a�9�v>�.E� ��>��B�p.7>��<�-����	>j�?��>q\?A2��j�>D�Ⱦ�:���e>�q5?0l�=��s?M�@?-��|�:��i>���>�*e������n���r�?$2�>�㭿�*3�@�?�甾�f�����ӏ�?���׋�>�`�=���>�ry���T={x?ٝ���`إ>Q��>�4i>�c���m>�"��h�=D�>�=��ۄ���$>{ �� ��L�������/��O��oO�XK�?�w]?��D?� >'K�Օc�v�J?�U��Q?[�_>�����>��?�l�>�4�>Y��>��>p_��4G�o��={�?��%?H$!>F��>?'}?��r��%���L��C�(=����R7I�d�?(~��>MIG��j4�Y5���>?�Uc�kF� �>��稾��ؾ�R@zs?��<�����{?��m���v���񾪆6@�;��3�<��|�?7|s�"`�Б)?�N>f�������Qн�4?`���9����h77>[�r�2Y>��&?;4��_��>���MD�K���?}��>=�~�Tpp�Z�J�.6�>�J��g�?j�4?��u>�h�>��=X�)��������t�=!�t>4f����?V��>�����#4�ٸ�?��i�n�5?�ߜ��(�V`?]x��o�þ��m�{�ǿ�O=��?6o���CȾ�\�?�O�Ԍ�M�L��">�$>��I���_��=Z��?	D)>�ء��F7?��>G?c�����=�)���Ž��V�����`�?�[>>ZB<�o���>?B?}��y1�J��?�i��ta?�S ����'ɕ?;aI?X�P?����J�V>� ����Kt��) ��-7>h��>�^�(Mw�Mq?]�\D�KN�>K�?��?*��>֝�>�W�?�(�>8i�>�F>������d����>&�>N�o?"|W>���=$Ͱ�`���!}�ه�m�9��҆��N�Em���'�� �{��o�?e��=��ӽ� ���C����ו�&�#?���J4�>�~�?�Y�?6�?��>K�h?i_����@?�K=>�T?O�Q���M?�r�:G_?n�?|�m�ܠ}>��a����Wn�f��?D��>�h?d���h,�?g��?�ܚ?���j��?���_9�n���k7?EԠ>�����M?��g�ۍ_?|BM=�(?��X=l?���l0����?٦?9{�>�����0"?�I(�O/h?�㩾͖̾�Dӿ�D?b�M�0�����h����?�i=���E=I�ۿ1Fx���C�2i�C]	�W��������=u����I�?�a}=��?�e�>��E?<I��e���Y`>��g?Y�O��|q>|�?�Y>�?i�?�e���H��W������K?խ<�)�?b��=�|����>AM?�c1?�ST�I_�>:5-?�y���V?���>y�%>!�K���a�m�j>/��?�nX?6�D������,z���H��=��*�_�S�&��?E����<�~�\?O]Z?�TZ>矕�a.?8Q?�N�>������?��> 
?I	��-?���iԾ�kϾZ�����о	읾A�"�	>;�?�P?�J�>pg�>4c�>w���t弮'$=�À�}c׾�C�>�P$=�E*�G��͍S���ݾ%�d??-�=2!�?�Z���8s?sݕ>�n�?��r�H���`��>N�����~?7q�>�A�?p7�>5j=���U<��q�ݾ�Ie?@p��8��=��?�g`?uפ?�,?�n׾V�>�m�?M�c?��ƻ�-�Ͼ���?f
�>�	��%~>�~��?��?�ƾ{�[�?-?x� ?�پ����\>�  ��d�>L�[=~�w��<�=?��?�Ry��?OT@j�׾��Z=��q��+�9�e�Z�&>�?�Ȱ?���?�R��.�1�?�D��I�e&�5�����>-��>�?�>���c�μ�'�R������>E�&?���͉徵��=YST?��?>!?O��?�h\?�� �
�=�5�>�'�?V�?�D*���??tA��BH����I��`jN?I�'>��U>��=E�V���r��&�=����l?/����x>/��>Qڞ��᪾�� �o�>�ev�Y������|?D�����|�Rɥ>�^?�쨾��*���.�O��>3b`����>ʥ?���>r�@�{�e�����a?�v;;�G�<��A�
ƭ?2�4�%�����N�.�?���> ?�?NQ3?�3y��d&>��?����]���>�G(?�N&��bP?�����m>(�ྙ4־�+<4M�U���>g?�?ժ�M��>@Z��&���Ҿר��� =S��=�^>��H?��׿##��L�0�,��ۜ?�o"?sK�?� ��F_�?��>�Ò�h`Ǿ�h ��R���u��(?�h2?B��?��^=�wz?��5>���"�)�@�!��(��o�>�,v?PCM?���>�۩>�¿��ƿ�آ?�p�>��U?q�#?�^�ӐL�ln>=�?���>k{?�6?�c? 3��^Ѭ=/&:>�<x�?��yW�4Ӟ������*���2q���K?���<�e$�zè>)k?�A�?:L}>�o���>�����b��ѩ5�g��?[�A�W����u_�1A?���;j}I��t��5�-�
_�<O*?1r�>��?r�S��-)�Lof�M�\.Z?�@F��?���?rh?ޱ?(��� �����)�=>�S�@L?�@���]�i0��eW4���?�q>��?�K������>�9>��>�>���?r]�?�ľC��7��e�>���fK^�rKӾ�v+��k���Ӷ=��?k���f��,�f�Ӣ�����Y^���i������j��y��S��e��?W�E��5l?F���AN?W
ÿ�P�<� ��=�@����.G�>��������x@��W	?�~��}?�?_�>�.?��@�} @�*�?�4�>��?��?�� ?�����?���>��M��?m*?��+�	+��_���9L�?A(ؿ��?���?W�>�i���S?��?W����?����L��>U����(?�*G�پ�?�>$L?$��t�=����>�x?��@U!
@>��?k�? �j>,d��G�#���&�)y�> wa�k����׾�9ѿe�? U�?��x�i�?�o-�5�;&)?�?a�i>��-�P�>G��>�Ⱦ>v?mF?�0��2�)�@=o?���=:˦?/._?�P?z!�j��e	?G��Q�?����?���s�>��	�q��?��̿?�>�wF�Ɏ_?����k.?4��>G�9��0:='�A?b���Z�B��f8?��?����n�$)���E����]���[��Z?��b>�d�@FD����>Q�>��>e��X�ھ�b��cb���>�޾>N �?������Q?)��C���b=ɍ&=m�߽�UV�٤e>*pȿ��?��J?�`�?}<,�^�7��?����N�6a�>Ջ�<�C?;!���W�>��>@�?]�>����#��IJ�>>�>d��?�ZY�6Ҿ���!�?�9����!��E�>�ȸ?�|r�cQ>
9�>��=���H�����)������z�P�\?�A�?L<K@�d4�?��?؏��� ̿}s���N��a�B�N;Lb?fR?�{c��K��Vn�[f��Ť������\��1Dl�r��>O
�?U�5?�?�N��B�=�v�> ���.�Z?��{?��3?)��=��d�4e!> E;����=5�2�zZ����>��>�M=��X�U�0��>VO�?���>��a?2�>c����>8�0��_��ߛS����hn��OE>�K1>*i�����A�<�;��$?��?Н�>�:?�‿��	?�z����=�K��E뻿$�>k�L��Ą=�a>Ce��SQT?�U�B�H��)?9�	�ϲ�iJ�>��?n��>�h�?qG��㵾t?q��>|	�?ے����*>%��U�>�9�=v	�T��o��E¤��;q7����w>p�?>
?XZ�>G��?q^i��"�>F�>fq>M~5?��b�*�>����쏩����>˷.��Lh?�=>@@a��r�>B]�ॢ��*N�O���!H�?�ל�̒�?��?��R�S����ZпuZ�?�zc��}?�J�=W��?2��?�q@>CM@[(�=�����ַ�=�#��r�� >�ދ�!Q�,�z�-=8�i�ȑ)�Z\¾�q!��P��=Tʰ��8 >K�>�_?�>���91?���j��>����_�2�c8��)�=�w8�b�����C�m������¾-�8����=�L]>�3�=
3�����=��=��1�3�:4R>�(>{�>�i�>]�>��6=*r�>l���x��x�=�!R?f��= ^��H�,>è+>f��>��6����C|=SDR�D]���J��l� ��}���tվ�ץ�r��=��{>j�?>%t��9�-=r�>�+k>ҏS�VVE?���W�>Md�>�U>����bO0>$��=f�������{�<�m>�ٔ�Ww����>i�=��?�S�t-6>���ѾO�����=l�;�� E>ӾͶL�;��=��W;�����i=f�>���>�K>>$��>�f龨m��I̒>ݱ�9l(����4�<�M�=������5��5�>�SL=KG��(U���־���>���>�Td>U�>�g#>4�5���43>�=q�l���ľWɓ=Ѥ>����=�������=`E=q��a]�]�>�Q��O�Ž):�K�f>=����[#>F����a>�_=�T0>%�=�Y�>0d�{�_=)C��F�� ���>y݆>��f�7�=�	=��>b-�w%����<�~n=�>�~~���{�0Ͼ�!Ͼ�~��h�>8#�=b\��D�S���]>B
>7.�jѥ>�b�|�>,V���R>��1?�_=�򹾆F�=%��>q�>�a��hǽ�Ѓ>�d��w��̝[��D9=�z�⼸����D���~�T����CB<T��>���=s�����>�U
?��?>��[`=�w3>p�c>(o��jK�>�=�>���>��$>��>���%��w�B�{��>�:��9��;`��CM>%���2.>W����mǼ����ί>�?�e��;� �G�>�3�>�m>����D3�=]��>^�>�nT=x��>�E?�6U>��=C:�>�q>����G辒�0>���>P^�	>��[�<j�>�>'<e�~W9�g)�>�x���E>rnN?���>{���o?��ǽ`c@?�ހ��GԻ�}��H?Ul3>����̮7���a�G��U�A��K���[�D��{�����6>����(����y=y��>��!>��Y�sJ?Ib���s�>� ?Y]:?ab�q"���I>���>���=vҋ�n�'�j^3=�Q[�+���������̾	�}�\����Ͻi�ʽ�	�>1@?i�`����>��P�y�G?���i@4�P�`�ס�>7��K�]���ݼ.��YQ>�&��*�=��>�빽����<�3�L>���܉���Q����>*$'<"h�=?޼=���>C��=��>�F�>C7>�=3���k�>��>�T��R�'�q����4>��ϽM+���Ӿ(����P>c咽%���PJ�>]�ƽq�þk���b�E>f8�<�����գW>sĊ=Ai���<>���>wp�<�#�$�ƾ\�;>(��m6>�ľ���=
*>�w��@�����=���>�0�>���>�%�>����������h(>�2�\<>����Q=iܻ=!NE=%�T�s=h�>�ۼ>�Į>��>�q>���Ce�!b>s���Ij��տ�S��=�f=�-����½Jc�>N>$�Q>TU>���>��=�6�>��u"����V>Ojv��\C����v.��v���U_��}쾿�j�8�[����*%�����V�پ�b��ɷe��Ia�H䡾�M�;lJ>��>�V��%�ƾ�s�b>˳s����̓�=�ة>R��>��*?�;����>��=5��&	����=�=�@r��+�J���
_�t�= =b>�v�>B��O��>�4���|�>L���>룽�׹=8�=�|��eƾ'Н��`d�O�����>W��=U�C��Ƣ��/�>�+��<���c���>�jh�D�T<WW(=� �>u�>��==r��>uY�>��=��W���=�gH>�@�����mt�+��>����|5�䧤<�j�>vh=��=���>򲎾��.��+�<� �>JbF=~��}e�|�>j+> �k��{Q=�.�>��>MJ�>�r�>���>�`p=\��>�v?#��y�E?�@�o[�>�Ո<�S�_K���1>e�=휾4�c��t<�cE7���=O��>���>K�f��S�>�1>73�>�M���>P^ܽ�Ӄ>S��=�ڣ<�8���>I�C�u��>܈����䛍>Ch¾���>]��s&Q>���>��?��;�(�=w��>x
X>�I�>�*?�;��1.�P��d�潻�C�D�o��y�����>�[>�s����p/�|�3>�5C����2L�KcZ�b[>��1?�=��	P>���E;��?�=�k��aH��o�>�_�=qʾ�	�W����>��̾pZ=؎\>t>�`��5��>ɝy�٫�>��w��<���<f<
��=q�žs�����O��{����=a?R�?V�����?N}���?�+>��<�,��N�>U�Y>��\�&/[>��G�2f��-K�>��?1�&��#���$�YV%?�B=�~�K���u�#>M��䳟��z���̽��V��d���*�>6$?+Ψ>��T?_�4?t�8?�C�>���>GvP?��u?�>Ol>�"�=JCE?|Ը>��>�~��*]�=��.?���>7��I�?��)��(D?�E���[=� 4��?�#��Y�����=s��>���W���3��巰�S�]�=�z>}�(����z�==Ok>>K$����Q�K�{<kMn<u�̾�=�z�>V�>�Ǿ#R�>{�>(��>�[ ���>%�6��i�>G���}.��9߂�w{��צ������۾	1����=[X��=I>O�1�񧀾��.>���=+Ҵ��_�n��==����:�yO>4�->���>�~e�^e��Q��=x~?��[>c܂�uO>)��>++=����D/��->�0��X��coƾ�����x��E�e2���Q�>�]�����0o��Y�1>�6>8JѾ���=]�<��7�
�о�H��v�9�?��>T�@>U0����@>�>/;�>���^ �>�sܽQj
?ު����=d����'�>�:]>S��[���l��>u_��M��x���2�>ď�8X>��-H> LB>��^>��<O��>ō��y/���? �?6z¾%?'�u��e?�]�51<��{���J�>	9,��=����U	��%`��лm �>�Q�>!2p�[�?S����	?�p'��d�v��m�~>�=r���c�8��3�'����=AǾ�{>�y�>#+.��/=��Ľ>-�>M�>1����M<%�5=�ֽ��=�e>�F2��O��d�B<���>{)8��j,>���>�[�>�!q>��>$�>�u�>)&>�[�>�!�>�C?��X?�OԽ�AA�306��J?��|>�(��U�U�?q>�:��%S�=J�׽3��D�¾4�۾�����Z�zf��PνTGK>��>�=��:�� >u>�Z�ȫ��OӢ�W�2>ͼ��<����(�޾��>n(4��Q>j%��?@/�-{>�H�=�;�NLQ<�g�>�cc>���>�>��d>�Ǌ>���=S�>B�P>àx����>V�+37>_)ǽI��~(��x�B=#���5�=����^�>I`?Γ���Θ�e�U���>�|�ᖀ�X��+I�=Y��PdD�bݙ�n�;��Gt����|���[��)矾��l�� >���> 51�����<� >5dN��u��&޼[t�<�%ؾ��I���/7�O'Z�!��>�x=>���>���jq>����r>�ܩ�kV�<�\����9>�[�>Jf�>���>���>�S>�q�Jܾ��v�'�>v���ҕv�\�����=��T���=N��D9�&"���z����^=�"�3��=�[f��>[���VU��6�#!�?�U���=�Ԍ���>h]Ѿ[���)C����?�A���ȿU�#@w/?�]��6>��>1�F���@.pJ��.��=q*��̪>+��>8�d?�@ҡ�?]�=���?�?.�Y?�C��Dy%?Wu�><$�����Y�?
 �W�ٿ�Z��<.����B��!�� ��>�Ϸ?������y�>���?�7 >W��?T2'>�̵���>���?6ee?�h�>��i�f灿Q�1?y�j�-��$��Sؾ��)���4>&�T�:���?Y���@[��ȥ��ֿ`"�c_>���?�|@ۊ��:?�[q����?S(����>Hiƾr����iG>RM;�h7?�A?�E9�n��h����*�<徾���=����4?s�H���1�u�1?��4?�?�럼�2���b���֎>�D?f�8�"�A�g]�>p�H�@�۽��?�U�?"݊?��m?_q��M꺿"Y?Ѣ�?��¾�����/�?��}>E	�����t�I���I����(W�z�>>�pt>�<>۩����j9������E�?�Y޿$��?k�>Dj�?�(�9���&�?��,3�<;)?<��>X?��>mu=<�����F>5w�?rǏ?�o�>���<�>9�N?�=�?m�]��dw>�翳/@>���{^?�c?������k�D�ci�MD�>"٭?�:%�-�-@o:ξ`D_?��;)�����3���=�^,>��?�A�>F����*E?��ҿҭ��C1?�}S���d?@ı>^U�r-���?	@E�5��a���k�3�?�Β��އ>���6d(?�@����?���!@_���)vھ���=�$�����ȿ�� �����1��?U�>��>��?��["����?Ѥ?�h�?>�?��D?ң�?���?t�C?��T?��̾vAտ_�y���>/{"?} s��	?�{?ڟ���6�����S^�7#�"�����?�zm?I���7�#�� �?(�@�$���2��F�?yܚ�����**?v9?&�?Ts�>	?#z?�Wſ����D����>"��>Hq޿'�M?����t��?�?5�?7��?&~��$y�?V�=v�>�b>�20P?!R=�Eབྷ�ܿ��?�Bk?hȳ�ϸ��P���xS>#\3�L� ��L�>A���n� ��`�?#޾ K=�}2�Әo?M�Q�Qx��F�?P"�p�>���s��n9�����"@�'�?@�?j&�?�(��g�>�q�;��=��=?�)?�2��k��To˾"�=p8�?=��>kRU>�<?�hB��ę=\��?a��?���?٥�=kp����?߫�?���=�ߑ?�̾��_?�;�>�\'>��t���ռ<�H?�ҿ
�W��N�>�&8?�%�'a$=
[��sS?��=I��?�2�<�e>B_?�܄?�z�?vy�@ȩ�5f��H�>@�	?��k�V=�>SΌ��Zv�P>�0E?���>��>�]�>E6����{�e꛾�����R?%���ye?�o?�i��Ą����3|9>.ǡ�x�?�д�	U	���>�kv?̳���Ҳ>�e������=n����0?q����?w��=��K>l�j?f���=��4�?����*���<7�??_^ſ��;?�$��3?%聿�y�=�Ў���G>���?��>����f�"�[����X�����i�>�����o}���{?���?V�m��=��,��2�?kx=f�=�(F���`��k����?60�?e�>@s;���?n?�;w?0i����/�e�Y��,�?M����@���G[!?v9	>��?P�?��p�����*�1>=�>?���"����þ�*�>i��?��?�(�?(B?1)����?K��>;e=?\z�%�۾�l�c��(�����c�>t@��J���?���?���S���x�>$u��΄>"��?��U�,�*����B���?�H�>V�Խ�~p>ߩ<>��1�����4�=V���۫����>t:�;<���V����ۼ�4�>��?��B=�u>᠛���/>8d��ޑ�N*=^��=	�޿=�>������E?�bS��j�iu�?'��=:�����?hڎ�X};?��m�N�
cJ�溋�Y�-���=�7�<����r;B����;ξ��yN0>R��?ә.?���?��?�7���> t�>��V?f�>v(���I?�����2��;/����>TmG��N�������v����?� �?j��>`�?�*�?Q�>��޾���>�� �%&žH-?c�@z�?���KR׾��(>���>�
?vZ^>>-{?d��?$�:|��?+S}>�Yx>�5;?�-?��+��%r���ǿ;�O>p�?d�?<=�?�0T���w���Ⱦ���ZD�>�B<?�Y�����B���ǂ�$��? D��*T�|A���ȿ?j�[>P�C>�&�����??z��Br�?�(�>ό�?#E`�������=�t�?��H�q�]?�9�>��?}��ҍ#���t5?�ȿ�|�=m&<?A >&��PL�?�f��H��>`����a>cyE��J���?�fR?Z��?�`���V��0�¿n˽M�\�aR>��?B֫���=��?:��?��>?�?׽��x?����-xɽ�	�ar?�?�2ת>�� �|p˾�G.>)k*��>���m�?R�k�7ܰ?!��Z�b>�r>_T���TӼ��?��d?�ؽl+����HɅ?z����(�?�Z��.[�?�Ӄ>�:`>{��%��=�b�>9�ÿ����􃾣/S>kp~������O	��(�> ����@Y�h��?�?��>��>�:�>�=?��W�4i�>�>�_">�Ǿ�6�Yqc���>���?U��~�9?#�&?ڇо�¾O�Y�p�?W�5��{��)����?�ݓ?�x�=�D���=t�¿��ο�/`�(��P~����¾b*"��v��V��?�P?F?��??��?�Q���=����?�9?>���U>_�?b�o>}�!�A�>�����>���l7N����>O"�>q����8�\(��1l>�HO<�n��V8
?;��=�K�u�
@r	`>2峾���?��$>�%?��P<Ə���(�&�>�2�?�鿳��?;*!���p=��d��]�?%�A>|�ֽ���#�>N�@���=�H���韾�bw?�1c?"k?eO��x௿F�=?���<W8����gJf?*�?l���?$ǖ>9�B�aD��+�>O�>~�>�ύ=��,�J�?3�>�Hv����=d��?䤬�=��[]�?6p;?s'����j�/gd<�����;?|+>��S�?^�?��n)?�a7?�"?������?)�l>�/S?�WR�v�?�h�����H��O*G���>4��=�v��a<�'�Z0�?MU>�Ӿ|L˼���+�@T��GP����?��ƿ	ە�A,?��?�hh?��;c綿z�l�`q��{;>P}E?RaN���&�x�?u�V=�S�ix?��=��>yִ�"�?C�?^7w�S�o���>��j��[2����y�-�9��cZ�7,�5�>uT�>��u?jӧ?��=Tl�=o��=!�?�[��V]s?$?��R�*H�>�m�yP�������C���j?/i�姾��w?4�ȿ���r�q?���>P�">��:$�����_G����=���~�];���?�26��L�j&���ѽuB���>վ���)�	?�X7��>���q@�iվ����׶?_ �����;���G�k?W�r>�v?�f��c���lE?Q\?��|j?�T,?�~ֿ��E�iD"?��"=�P.?Ơ.�. 	�
{m?fp�={2�?��+�Ž��ݾb#�>U?ʾ��c���=Kp1��� �9��pp<@Ht ?3y����B.�����?�ƿ��97�L>�e->���>�Uw?�3>,�ྻ����C>�ԾgA?P|�?�?��>��1����PL�?ߚ��e|�?u��?��&>��>�����?TSD�*��>�P��O@5ſ��x?8��?K�\>8����]�>PK&{�<      PK                      archive/data/8FB  á,��^�y^��!_���+�<��1������@�������������(��M��>�(�a���j>or��S}Y��q)�PN��
�|�Mo��6R���|�g>���
���ؾ���]�e��5�2����E���K��~L�U��0C�z��a����>�25��M�:T/����m�>�|��d�)�!a����������֥2�b⡼��2�EJ����?2�$���D��-�׾�S��O?�阿�R�_��vr�������f{ �a����4��wQ����6�2�����R˔��������]�''Q�a��1 �" ?�(�A��>����y��\��98��%�=�|���0���-��,���P���߾�ľ2�"V�>�-�?�B���C�@���`����Q�g_?�9��0���Ho>ϟ*��"��\L�A�_M�X�>�����x!�<6U�r�k��ds���"�������1��x��}�>:���}�PKey�O      PK                      archive/data/9FB  <Aͽ�@��&�e=��l>�I4��_>α,�9 ཎ}>I<�K���)>��>�hC>�[�>��?�v��xF>*˻�����o<�G�=�¡>^�>���=k�>�?��k;0u?2�>��@�=.Q?q)�>OR��\���>B��iI��-<?7��=3�`<u=?j�>>�4>-M�>"�:+ �>o��>Մ����<
�}����:�="^>�a,�e�>���>�<b�˽4�:F�F���>w{�Vp�>�ê<j�4>"��<���;�_K=G�D?�u��G��e/<6���c�>�-�4g}=�8��l�E <�����<J�?B��=�ݱ>#_�P���|��=c�c>9�?�`��P&?�}�=ĩ^��$9��NS��r�=���>�M5?[��>��σ���7�>y~?Ǳ[����=��?��-�)��>cL�=�;?���>&��>�C�����>C�I>o�>�I>��==;�=��ʾt)z=[:#?��@����=x�Ľ���
D�+EP��������=����1'��==�d��1��>*O�>p�	�񁇽��+>���>d�=0/�>���>YI���N>G��%8�>�ˁ�r�W>�>�>�r>�f��$�>�x��=��9��U�>��<��g��a�=�\�=~���M>�{ ?��<��s>Ʈ>Yr����>�z�>�����?���:ƪv>-�R>�Q����=��>w2'>�*? e?���>:5?=��=���>�G�<)M�>I~�>C��u�>�<���>��<��9��1<��=�c�=7O*��.v<��>�2��9��<��ɾ��꽅�x�.f2<u7 =r�=�ߡ>5N ?�B����������>.�_=p�?�p�>r�=p�1>fx<�Y=�>iݾ;��?�X��o?r>>�����0�餽c�V?�a�=g"�>S{���!Q���>�6��-�E?ڮ��5<�x/?�k�>���>���>�<��Ճ>�%��ws�-�=��?�w!?���>V������>]"�P���������>~��>�-
��dy?�ey�je�<�S�>�fm> Z��}�>*?�&=?	*�?4?��ǽ�>x�8��MM>uR�:�p�zu?�s�D���]a<���>_,����=*�n>?m���M��B*>���>m�"��T?q���ĸ��>_u�={Y�>���>��>~(�>�_?�]����>�־>��r?��2=��I�1�?aþ�=G�?��>��	?�?�<�4ؾ:5����=��=��U��h�>�q<&}�>pqʺ�p� ���W��naD���?��~,;d}j��Q�������"��$�>l�>H�뽜pD=�k�<�L�>%?�p?& ������?��>�)�>�ۭ>�Kļ����͒>>5g�>&�ۼ��>u��3�8?�s�I�H?���>��>��j>�~�>��>I�X�$�����>��=��R?�.�z�����>��>���>#h�=�G�Nh?6�%�p�>(Q<�G^=�A-?���>�9�=x�?�֬����=�樾�坾���zW�"���;�r>Nw*��[�>l��>��	?��!?LP�>�\���>���>Zj���o���o=Fp�>ia@=F[>Z����8&=�c�ph�c�>|��<ߟ龌�A?�r$<@�+�e���x�>SH��]
?oΟ>��<(�N��2>ܼ���? d�>zBD?q?��=5mａ�־>H>�G�c�z=�������>���a �r��>�3?ZE~<E�g��<����s�>�G��W���M���o�>Enz�gPּ3�>֣M>&T�>�g�>��H�[! >D��=�%�����_���S)>���>[4�y��<�c?��Ͻ:K=������>9�߽�s����	:��E�Ay:x�>���<
e�?�e?o��M�=?L�J���k>�=t��>�6?�P�>4�O!�����>?W?�6�>,�A>��0���S�X �>��>�¹�����D�!��<�y�>2�b��;��2�N>`�>���==�PKL�      PK                     C archive/versionFB? ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ3
PKўgU      PK          ����                     archive/data.pklPK          4'f �   �               R  archive/data/0PK          ��Yd                   Д  archive/data/1PK          ����                   �  archive/data/10PK          
��2                   ��  archive/data/2PK          Y��                   �  archive/data/3PK          ��c4                   P�  archive/data/4PK          [o;                   ��  archive/data/5PK          Ƶ��                   Л  archive/data/6PK          &{�<                   �  archive/data/7PK          ey�O                   �� archive/data/8PK          L�                   О archive/data/9PK          ўgU                   � archive/versionPK,       -                             ��     PK    ��        PK        ��   