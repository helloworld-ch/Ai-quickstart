PK                      archive/data.pklFB ZZZZZZZZZZZZZZ�ccollections
OrderedDict
q )Rq(X
   fc1.weightqctorch._utils
_rebuild_tensor_v2
q((X   storageqctorch
FloatStorage
qX   0qX   cpuqM tqQK K@K�q	KK�q
�h )RqtqRqX   fc1.biasqh((hhX   1qhK@tqQK K@�qK�q�h )RqtqRqX
   fc2.weightqh((hhX   2qhM  tqQK K�K@�qK@K�q�h )RqtqRqX   fc2.biasqh((hhX   3qhK�tq QK K��q!K�q"�h )Rq#tq$Rq%X
   out.weightq&h((hhX   4q'hM tq(QK KK��q)K�K�q*�h )Rq+tq,Rq-X   out.biasq.h((hhX   5q/hKtq0QK K�q1K�q2�h )Rq3tq4Rq5u}q6X	   _metadataq7h )Rq8(X    q9}q:X   versionq;KsX   fc1q<}q=h;KsX   fc2q>}q?h;KsX   outq@}qAh;Ksusb.PK�od�p  p  PK                      archive/data/0FB ZZZZZZZZZZZZZZZZS�'��޻���\�$Y8���]�Q����#̿�p��S�4E���:�^8��[���Z�>��.>�����H?�(5@�� Ae�@/�/��$�@�D\@OF�@xN�@��d?;�l@� #����?%��@i,D�i��?�I$?�)��t+>��=1ޣ��$�o9�CL��G�/����;[���
��9v��7/�Z:�>����a�$V��"�$��0 �1��5�b>�xt���1>��ʽ�� �;DǾX����Q>cC˾�ף=E�2���%�R����އ�W3�F߿�&?�-;��3��mt\>�)��E+>xnw>:(&��v���L>��Ƽ��=�:�=�	��(MJ�ޜM>Nv����0=~(�������>^QX�扭=�T�!�>�i,���h@�@�V"@�OS@�^�@�ђ@�£@)$�@�м?S�W@x�@�J�@�@�X�@�.�@2�a@#w@��@���?r��*�@u�K@�(8=��@?-�@ʁ���gM?�y��L��ٴ�;m�?�30�.�K����'r�����g��=��)�_�.}��
t۽�B���B?�\D�e�v>�����I��J������U����(�>�W迀L;�w���\��"X�'@��b��f�V���e����Ly�T��Jzӿ�U$�L'ҿサ�T�>��P�r���b&���O�*���B����*?(��������B��ٕV������4��n����qJ�(g��\�Q���>�bu=jH�����<��EL��O�[�K�y`�=V�<>�t��T?��@4�;@�;X?�wi��^L��$�>4�L���م� �B�y�ҿ�6����?����ت>w�H@s�]�������?�*��D��;��<̿_���T��H���^n�?q�#?t�п�.k>�L@~@Ƣ)@kA��?Y[�@�G3���@���,�9@�3{��ۮ?��@6l9@�@厮����?�)���ҿJ�i�A�Y���<��t��87�ߨ���>b���A��U�W�O�����?����n�:�����>�B���L
�~�����0�<���%�6�L�:��>�z�XJ��O6��Z�� Y>� /����@/�@�:��8�@���?��~��C @]>��=�f(Ͽ/F�7���$�?yq?���>ǽN?�Z?��Ϳd�@�y�?�b���p���5ŽW>H�QO�
^Q� ��I�p��@U�K�d�0o���@��}��\��O�����#�����b� ��n���ٰ��!����=`�r�:�������'�T߿@���:ſt9�>:�.?���kx>�驾��׿XAƿ`��� ���۾���>11h��~����>���������E=���3�L��$�CD��t]��p�=�O�CRj=.�>��|�9U���j1?+�Y@��>�2��mC)>?�L�B��?oJ��:x��3�?���?A.�@	'�?u(쿕2�?6��Iۿ���=u�b�.��۷)����jm2�G �E~t��TG���<���ۻ�����*�?��#��P�>�}��S"������Z���,�p�����\@��Q�Sf��T���Q��.^��T�5?� $�U��E���a��a*b���@J�0����?�`��JVG?���>�F�?��x@��?��侳y�?	?�@�@|,�?��+���鼼Լ��?� 	9�?���A2ᾠ�}?K�?���:�ٿ�>ľL6��%?<�&����Cd?�Tþ����3��J��nx=�J�M����h/�=�����ʱ��^Q��F�쐵�i
?ͦ�@l��@}�@��@dU)@��j@��p@�L�@�#
@P�Al�@�58@�]@� @�87@�t�?��@��?�Q
>U��?1�ӿi�Gv��]Ws@������?k��?_�F���ο�UV�����E�*��r���J������D>��A>@����}� v��� gּx�;�P+���=P�R�Č���/@�� @�!A��4@C�@�W��ɧ@�u4���)@�V3@K��?T��=�W|?D)�@{0�@���?�䯿y�Y�J�q�Dvھ�7o���>��1�Q�%����-a�}�
?&�=i៿��/�=�`�(zz� �4�)o=ܳԽ ]=��=���;�(=���=a�9�s%���e=�ƌ=t�7>>�߽�b#�+�!@ ����k?n���7����Y&?覠>%��?�K�?ҧ�2U��`E�uUu?�l,@�O�.k�>-�V@��@�"������G@���@j��d�?�8�@-�@ᕛ?�$�?���@���@�@��A�^C��FQ=M3L>�n��t���<Bs]�|F�=���=0�Ӽ��E��&��b=�Ke�x�l�`PS���B���H�yh�l�<�U޽�=��'�E�=�V<� �e4=�~=���-u����\��(�.�S>�'"���9���b�{]��V��Ѩ��|@��y�&���J��v��� �a���t>��>��S?������������^��,���IE��l��!��y����o����"J�t,���q����I�ٿx2�����)S�!�2�(��;,����?p��R��9������K���06�?ao?S�M��7V��t��[��d�>!0��?��<���BR�x#�#EG���˿�D��4��[���ih������b@	@9U=�4r@
�@�q�@.v�@����^�@Ұ�@�}�@��g�:@��(�?���@s��ƻ�4��g�M���n��{��W�d�q�����	�}��j> ?.C�>�᭾�n����?�
b@�>�?|�7@�؟@�s�M��?y@T�W@U`���]V��*@::�?���?_��@�#���ɧ@��@���@a�p�lV@!�@�`ɿZ�� )@%����6ƿ��?Eƃ�	��?L�?�	;@x�\�/�=��=Yǹ���2�L7����=�8�=;QL=(A��f^=����n��z(A>��<��Z��R@3c|@'ur?���?aQ�?:�t?�nĿ�~k��3z�0T	=~�����@��u��m�?$��@Y��@���>n��vC��C{n����B�E����������/i�W�4��̿��5��n:�c��rlG���@��e?l���]��D�ȹȢZ�k��?�D?�)�q���^��p�@ݑT��2����6���?��@9
@��H�R��?��|?{3->ގ�?2�C@\k�b���k����E?�q ��~�@���>T�k���@L�?��R������@�X@�6�@�ٙ�8�4��f�?�[@������?��9@�O@itܾ.��>�_�>�&���?��<s��?�����x�?���V̔?��A�:?�\'?��l��O��'��=��f�F^�=(Q��z�=?Z��i�ѽ�*>���?.M=7��=�����w{���=̻��Xxz�(=��)=8�n��:y��@� h���=����<����"�<���>a=`7����^\�=3���CD�������I�q��V�y�x��=Z��:OF�σ�=�>���E3�>#Cؿ�e���=���>��G�}�3��� ��B�D�O�,"��48�>� ?mJ?��C?�j�p+J�����ӾG�?-�&�h�*�`ϟ>�誽T =�W��˲���6��2~����ۿN��>	�
HZ>c޹�����;e>�uW�3c���,���5�D���u���[e�w����?�*[��������;���A�<-:5������sꏽ��?X�!?Ӥ�6ʞ�A�)��)X��?W��Dk?�&�?S]g�#���@��o��Cq�?J�C�(W����=J�W�f!�sY��>�0rӽ�k�=��Z��,f���:��h���K��`���̽h�&?F&�Np/�V&����?���>�d署M�	N�>��翐��?^v�? �>�.�Z#;X����<e>�cx?>��>�-@�(��]Qʾ	��?��@�.�/�,ϖ�)(@���?h��<�-
��1����=�$=]P����=>���0����(+3���C��b�>YL���l�U������� �gG?PK�O#�      PK                      archive/data/1FB  ��
���M��.������o߾�q��J���gҨ���<���+?���������b��@�ӏ��������@ѹ�@��@�ꝾE� �F��GG��)@�����;��Y��x��̯�@D�X���,���O��^��-��@������S�[r��U���;�@m�L�C�ŽU8q�I\]�O�ǿ*}��Â���@C?:�Ͽ:�@��l�ȣ��P�@e���E�o
#�w�T�b��@��⾒E����ͽ�@�yr�PK����      PK                      archive/data/2FB  3<�>Iܔ?1�=��8(�<N꽩4ɿ��ҿ��=�{¾ȭ=Б�5ٟ���?\L��6��)��L>�o���?�J��N��=K���r?�b�>�%W=�|=���s����c_�ċ�=yϒ��3�=���=��8��f���ӽ*��"���Q��q�b?�2!��p��`�/�ϑ7@�Kc���ν@e�?s�?6�?���?��9=X$�=x(#=5�z�\&�=�θ=b6���a�;��=��'����/e�=I�?ym�?W� Ň��Ӫ��oͽ� ����?
?���
Ŀ�,=r �>�{>7���&�,�?�оѦN��J>-l�?>G&����ْ��e�>�վ9|��{d?'l<GJ����RC��'Ŀiˑ? g� *ƿސǽ��=��5;�=$�>탿��>-�ؿ�*�60����L>d=k���{ ��%�>������>�^D?�<��p���>�R?�m;�%tv>H���b��yқ?��>�6q=0�j�Ԧ���>%� �.��=����y�B�� ����<��>l�>-J����c��{����_�����7�a6X=���[��`4����=�[��Y�=��X��K��'�<��a>Oj@�mF���U���C��z�4��=������=�bF=t+=,n�>דX�������������W�>��̽�<{=� ?i>2������XA �^}w�(������Bz�KR?��=y�;������<��@�aK�;^?X.ռǕ����=�T�����z^�=�ۊ�[�<�e��V��=��<|��S�A= ���C��=!�j�+)��\%��֡�� �=2+׽ �ͼ:��� �zd�� ]\:�U��,��9�������5��M���Gz�0}�=e�<S=����=�SP=U�=�=D��^���f�`��l_�C}5= �K���:��
���k<��E����p�G���=~`�={%�<������g�x�����=`����2Ƚبۼ��=���*������r��@��<O��J��<`�=��=��8���ҽ�������>�M:��4{�;쀓�B�� ���置��=)�[�<@�e�L=��½��º0�<�߽B�,���Y21��ߣ;�yۼB������½��r�f(�=T	��:�(�ndl=
&��y�����`=�%�=oϐ�&���h%�r�<��E�z��:�s�=,�N=*��`��{o����=OϽ[��<WŽ��ϽH��=�##�)������8â<�%��B6#�����q ��+�=a*������Z ={��u0�#��b�w�=���<�\�J:ϼT����!Y�՚�9R�	���5�f��<~[�0�:��KQ=�{	<f�=M?;�@}�;���=�޳�a~r��=�<H%�	,������QA��Հ�m;�=���=9�U=.���<�������V����^$�=(9��N&��ټ�Ž1@����e�|�-=��Ž0m<ԤƿN�-K|������7����{=Wۻ�`[�>&��=Cl����� �*���v>_]�?,@پ�H&���e��d���[�>,N:�А��F��= ��=[>�������ϡ�a�(=1Bپ���S�<�]�2.���� �Ճ�E���Y �8��<G_�FS�>kt.��IW���&��:�[�����>l��==FܿvL���z��U�V����)��.����}=����g�>ӡ<��K���]=��2=��*?����W�=9��?.��?6C�t=B���^��H�Q��?�ߧ;^G�?8�=v^�?�q>_�C�J?\ʘ��=~W�����=ُ��|A?�/t=��j��~b?���@>�Fi�W�Z���N>���=\��U{�T�4�(�v'h?$�-=��P;��G�$�I�� >c "�r.������g����m���=5���s{?��>���-?ľ�a�=���=��׾3[Q���{H�� $߼��<�t��(��4;�����>���?�?��#��l?���>�L�?���?ӂ!?���?����o�3�K��R�6�?J֕=���j�;��bm�>��M=�|���>>�Ǐ�Q����?����"Bs�4aV> ���2��������<z� ���@�(�_����f�ý��D=�у>��>Sw����>u��74:>�<hھ��H>�c?KY�ҼB?xo��Թսo�<�Ԑ�G�?�I?4M>��=�=W;P�ۚ���Z�>�Ʉ�A�@[��>1���	��=4ؼT{���)>�!�<��ڿ���> ��=7��¨�?*7[��=������g��}�ƾ��C?��?'��<������<(.��Q����������Q��\� 1��L�����Mx�=�<l��t�<���=�蟽&F�>]�?\��?Z3���x�'
I�6Q�+�>�}=8�࿿O�>+z�?"𫿱����������!=}�?��a?��=�y�(5.��{���� @(�e�W
=��j=�V�;�� ���3=�S�=��=^��{���:�=Gl�<��;vP��nׅ<��=$�m=Z�ƽЍ�<Ќ��=�����Z�<	�罠\���ǼL�ս�'%��K���[]���Ž 5;�X���Ľ�<�=%'"��C��Y�= �齈��<�����~C�С齘 x=��Q���� �=�8���ս.��G�<OK�2'L��tL�@��=Vs�=6L���oý�F�=�����~�= ��;��<گO���= &/<"��=���<_�Z<�<pڢ��,�ԗ��a�<k��= �����A���M����Z�	0�<��ֽ��}��<14�=C*g�`.#<��=<Խ�5��`=F�	��4�=�y����<؎�=���6�Ժ@f��:�����n��泽��ý��-��;�'�{�	�v�i�[��"i�= �;_K9=Xc�=0�����<���ύ��@�/��"ʽ�4�z���j/�1�<��ʼ�jg�ػl=k�Y�,���8!��\Ծ W�?�?�Q��⬽Z�j�_��J.�?B�>|h�?���oS���ʼ�����湾�/T�\��P�>Ν�?����l�
�������J>Bx0��6> ��>����K���Y��������jj(�F����2��X�; |��{�)��P?A�<�C6�� >�o|�͗���`c�8_6������>�fh��$�>�yh�(G�>Ӓ���0���=2W�=Y��?kn�>\����=`�j�fb���]�x�9?�90�L�>񽆾������>�Ǡ=����@�C=�?B	뽜�R?`>��x��?��@dy�A�����r,�����M�?�����ʞ>�w@�����>h��?�1��^E�0v��=����S� m=�3����F�,�p��=D9�<P��>C��'��>G:�>es>���?�	���=V+ÿ�g)����?����
wǿ ���ԃҽ$�=yˬ���?`₻Y2W?$�9��o�<���4_��_�=9�$?;��<�J]?�PA>@��=�R�<;�ƾ� d�ʐ?����?knW�2������ԿU�ѿ�-g=Q���.s�>�g��"s�>�n>9-�>zk����@?rt>�ݫ�?�@�>�K���??����a���:��~h�q
ͽ�賾,��=��x<V�����<��v��>�*��˛I?�Y��'}=\d��p#�}%�?�L�n4�m�)?�� �
��=��#���?���>/H�>�a�>μ�=��;�*���؞>KH�?�\��5ܿ��?ȧ$?�W;����)�x�zԾ6Z�?�V0?�L�?i,��P�(�}ü��`���>^��=T�ʾH>J)�>����L�/>.~�>b��)|E��@����B>-ڊ=wB��HR�=��
<}q�������<��>`����������=�^>)ы�?��<����>J��,=d�e��I�=�{��r�>���>VP���>��?�ƪ�y�={y�0&?��	)=n*���
=kʾ���?��r��>P?*�??�>W�?+��;��?�)?�?�?��ȿϾ�?g��#k���A���n#����?���>�ƞ��J�=�R�axG@]�V�%��>ؔ�?�g"�(1?������Cپy�?�W�>�bc=݈ѿȲ7�V`���)��=;��~��[����Y�99����R�st�?c�I�1��?�2�'�����=��=�#�>�n ?U(���п @�N¼e��<�̘�]�@�?�O?��<�$ޥ�I`�<b�\���Y?+�<���/�<�s�X
t=�֘��	�/w=��l������0�<�W���� ����lmG<=��<���S	��߼�
�0V(<��;ʢ�<�����2|��x#��O�<��ҽ�q�<�GM=0�<N�=�Y= p�8~�q=.=|�����3��:ء=��<������<΄Խ�z�<B�'��B�;X�м+	��H����C=Y��<��`;�e0����h��<���B�<Ab8����}B�=��?�d�����>�t�=+d���l�+O>g��?tS�6k�?�d���F߾np;�� ����M>�oO>��5��H����y����?Q�R>1�M�qs_?�L���2��1�`?->�5پI-��Hp4��j��5��k�=�UɽP��:D>�8<VW�??%��>�?���	:�=���b�i�K�b�`�S��W�>o�?4�Ǿ��&P��s=�(�=R`i?G�
@��>�c ?$�r�Ƚ�<�}[��"�?u�4��/��|��L^�d@{=�z=��ڿ�l>��F���W��|�=X�Ƚ����g����V�#�>�2�ʷ9�VJQ� ���� ���<�[Ƚ�$�=tƿ��!=�ɽM�˻��"�v;�?tt�a�?جt=h��<�`%����9J=B����6j���?Sq�����ɍ2�'���+ʿ���S=�4�>�CW?�I=��4�6s����B>8q-�0����Y=�fv���=b��?<=�8={J��@C�aCĽhG�<���=ʬ�=�>�=@��=��=7���r�<Ѿ���t���$��4=X޼:X@���Q�Ai�=��N�XK������~=y4��l=?K������豽�ͻ:��=8�i=2����<3=Xe��/ｰa�<���N��ѿ=
��Ɵ�=^)�;��𽑊��RZ==�y��=�����㼌�=�G=�ƽP�ֽQ���ŏ�/���xׯ=d�:=]����̼O���"�Ľ�n�
=�ͷ=���X�!���sx ��?�?�z�?���=��ۿ.�??.��?�.?3h�?TG?��n�b\9���l>����:־���g?ob�>倥�}�!>�����/ž79?:jQ?S�E�|$|�_v�>#f�;������/��=7Q��'*;��=���z&?y��=��|�*
н"��(�|>�k?�A����Ӽqk����<���>�걿�'��"G>(��=���=G�?�ZZ?�
�>	��T�� G<;���
y�>�(m?����Vɠ>��>��ڽY�>X�ｙ��<kW�?'F����`�}�\����f<�L�;7�Ƚ��?���=�7M?���Bȿ'T=�N�=Zj�>>�?P2R>0{�=����<Ϳ���x�۽����,�>TN�%0&?/�H������=�/>>�����5@�[��>�x��܈�<x�>�Z�>�;�=��4��܈����?�^F����=�?�+�h�ѽ�w �����ȧ�=ۡ�>�#�=����e�?���+�=m�^?�V;�I��K5�34;�NN�<�V>��|��>��?r~_?����K�n��}��-�>2%^��Ԫ�� �n-���Y>������>�5����cv�>�ס='�z��?};��E6���=Y��	}��A���v�y�[�_=x�����[?ۤ��14׿�g���M5�L�V��&?�ձ>���V1��v>���>0��п��ž�ŽJ���/?��Y?�;���$o>ph轤����=���	?H�]=�Z�=�ۼ�;i=0�Ļ'�n<"7�=�8��Z���Ax>x���%1&����=�?����@�����o>�i�AWb@0�@	�
@�oǽ���=wV���<���@}��K�����8���O�@~ͅ���$����<D�P=0��@,����S���|�<�T�>���@3��?�S�~��	@��%s��6���0��j!�@k��)��[@�4�������m=R&<UO���ƚ;͆=׃@�ȿm���?c��hl@�x��oϵ�Yi1� �����87�=�U�.�ɿ���ǣƽG^\�_L<��Ͻ~̅>�7�wA�Q�W�%n���C&�y>���<��;�F�=0E��=�
�_�0=��=��Խ��ݾO����ѽ�0��n��=>�̽R3��Y��@͕<���=���%�����	�����E���Q���yԢ>v4��@C��T�NvZ>�~�
�������@4���'����<56�<��>�֯=|�@=��N���=¦ >���>-�'?]$?M��> ❼K��=�6����H��:>��_�>�ƾ{;��'1ݾ]�־��X�����_#��b��>z�%���v?�&�=6Ǖ>�� �ٌ:>o�h=9����r>#x�>��/�4�1��|l�@���w~��>`N��ҖM��m�= B�;�W�>-?Խ��ž(�����>���>AD�>J�ͽ�	�:�?r��>gB�=)������0�>�3=cP=�)>1�
?����b>����B�=�9�=�����47��=d�:��cW��S��Fś=�p=|A��s����߽�Ɗ="_�=�:�nO��M=T�8=�4��x��t���н�%������<����Z?}�����J�*��=NU��L����׽,J�����2�=�t�hY콌�ֽ¼��н���,��=X8Լq~Ͻ�U��,ݽ�.=d�=�ዽȄ=�Tw<Z
���7���Wn=�K��4�����=Ky��G��;-���= bӼ;��AH��}4�㊉>Zܾ�<�����'��h<��� 9�<2l�(��?Q��<&u�w�����?��vɿ/D�B���u�<��T��3���a�<;�z?�R\�	�~?uB̿Վ?A�����B��z2?�h���r��Rƽ̧��)�?��>��= `�;g{K�omf<��[���p?��a�G�E? e.�C���
숽��ʿu`?Or?����O�>A`K?8�~=�B�=�^`=�U^>������S����=�E���#\?9�'�(���[>����?Ka��a�>r��?R)t���߿%f�?��?u^�����?����ۿ�5�=�T�׈�>c�'�=�;��#��V@vS2=�X���-?q!����b
뿬�x���v �����oh�00@���p��+��>�
�å=!��N� ?&$���н>�ܟ�i�J>em��~|�	V=�	���c�ޞ4�Î��@����ֿ秩=l����]��[�@Oo?��P��w��t���L�%N�>�?�ܐ�չ��xK>�7=����	=�ȿ.\�<i/�=�?}�*?�p7��Í��>�By�����=�@��a7@���<��@�?Q�F?<9�>˲=4�>��i=-ʿZD(?�X?��y�E'�J������QR�rýH$<���<z�=o��8�,?���֡����h�K�6>�,��q=�;�<�Z	��WN?[;,�H! �%(:?�!?�Y�������&?�_U?�g|����>��=���=��?��L�4��?q�佦y?��ӽ�t=xd�<�=|�=>�w�>��=�*�~��:�V����?�7о�sοS�?�ƽ:Co��G ?���{��������þܐ�=֨�_���J3���9�秿����㣽��ݽ�L�=��=�������߽�ʢ={]�=[A�ɸ�?�Oֽf����U>�Ͽ�_@Nx���j��U��_;�,���KT0��č� ���x�<����������$sY���2=>|A�;�����=
M�>��i���,��뵽^��<fR��G��(��s��>�MĽI��?_B�>�Jw��]?��
�{�-�4������[Ž��-?BO�?
�>
���6V�p-->oG)?�Ԑ� H������x�>�Q��O쬿"r��a�=���m=B��=P9$��k��eh�>>�ؾ.Z��V#>���{zK?���=ۄ=�9>�p��H�<?$���t?(Ɯ�ob��Tw=/}W?�av?!?�����P��
ޏ��E�=�>�g��mֿ]�=�s�U��j|𽁴�� 0)�E塽ǆ*?ZJ�9�N����������0? T=��>}�F���
>�:?ǽ ��F��^?��˽�4�#6����?�wa=�X�ۜ_��+|<�߽���vZ��n��>G�(a�=Z;�x��~?���'ؾP&����>���H��s���8�>=L6>��؁�?j�c�&�?���>�왽�р��ʚ�M�+��) ���r.۽0dü�|�5I|�)�U<��C��U�I��>D�>�=+���4舿z�<�n�)�u��?Ł>/��
�l>��	�$��=�b�>�U����	?�z?�����*�U�=҆��e�;�of�>^!�[�O���^� )ɽ!]O���Ѿ�>G5�<��m���=����彇9{�����O���=�Q�=�9�� X�8o�=��'>6�J���k�����?��s��q��pE�ܣ'�D?�b��d�8��z��=h��`6��{?�f=��̾�h�>��8?����}���B��f����?���>��?2Gt�u���*����������������.�L�>2>�?���=�s��%��ƾd=�Z���=	ͺ�侐m)����="$ҿۚ̿��=̲��F��=p`U�D膽��f?�sB��c>쾺<�ꭾ�7���"}=	9��n��K�?q,b>��>�
��~=��ҽX��<��V�����;��?*�0?�-ý  �b�E$A�[�ޝ?�ϴ���@9��?�Q7?�U?��L&�����ш8�h8�?:��?}�?)9��H�,���>��>�$c?Ę�2��ߟ!?�Q�Ro\��'l>�M>�@�?L�d�U�'�?kW?v���
�=z4���V��c���>R�<��>���V�0�����>�:=�S/Ŀo�*���?�/?�*�>�e����>p,�=�P�ċX>�ej��D1� �Pٹ��k�=ݏ<jUa�wټ?@E
��a�`��x��<��>먭�q�?�ur��v
�J�<�ܩ<��,=�5�=��ؿ����=*@�)�Ĕ=QH�?ؗ�?EcP��7+@9�X�QH��T�T�b8���m�:Gj�=�)9?l�5��j׾I�M�Q�?7]&�o䕿V�,�P��L-r����f�ͬ�?�>�>d%�=dou��0���@���>�f��)>йO>�3x�8 2��C��������=�(�?�	�������)׿�ڿ=�ɪ=���=�
�>�������l=�@��Mz�h��	�>=�Wʿ�֯��ˤ���?$D��o���r!8��FN����?��Z>�O@?����P�R��>U3�DA>;���咁��~ھ�vG? �s>�	���	�;�wy�h��?��s�--���z���ڿނ��>��=�W��~�(��f>C����H��쌽R�)<���>x(�>���Iԕ=�?�k=&Ї�H��ߤ�����>e�>��>?|D���>s�{�3�'��O��y��>��?a\'�Pˍ>`��;@
$��t�>������e?N� �,���2��=n����s�<�9�H��b���q�>�������=�j�?�,5,��<2�<
%׽�B���	>S�X�w�佻�O� ף�o�<=!���������=)b��	�:<�I=��X<�Lֽ@M~�nAr�4Xq= Z��`�Z���g=	M��l�^�ּ[�s���K<���<��<���=4\�ĝҽ�zT=\�_�Ko7�F���P͏�����Y�=��h½��!����=����Ҍ��&x=#���Fￓ�4�4|�?I5,?xs�>�S�=	���� �܄�?8�I?���?�ؼ���>4���|d��<?�����r��`���k?�E-?o����G�kM�?�I>��$�t��>�lS��uM� F�B]�=P�0��F���S<=8j��).�=���=3!=ur�>��3�3�u��f����>�>+���DY��� ��4|��4ph=�����W`�w�B<�`.�$��< DB�>[6?W[�?fM?�f>��R�t������h���?���J5><2[�;���<KX=���=�`���/���*=w��<��E��k0��=���0ŽNS)�n�q<�﬽)�V�z�)=^,=E�p��b��s��x O=�=�c]�c�j�=�%�0$���'�b��� ?q��IH����rŶ��k�=����.���6�j�=9q�n�Že���`=p1C��_��$�<�!�=��<a�t=���$2��y=�� �	�����;�	�;P��<F:Ľ�ؽb�2�+��=������?P�A?G@?��3?�B½��1���|?�F�?��>��y?ƇJ�o�.����f3�w��?�����Y��>�Qi�b @*�/=z��ho?l���^��CR�>���>OO�� ?��&�������*Ϳ����M�����}Q�=�b>஼�˾����,WD>9����5?�M��Sݼ�	н
��|�<�*�?�ӄ�C�>�;�� �=�A�������,�?Y�?7?0�R<`>��g���=���?b?�
����� ?KF=L���C�W��X���D��Y��Z���P7>j%��켿p�-�Dκ����3��=�p�rΘ�g�?�V������K�=��?��>���6ぽ\n�>�n��Z����k߽UB|�s��%\�;Y�h��<㒽|��̀�>�3>{~�=" �P�M�>��ݾ�8�=L�k=Z��>~�>H���4���xh��֮�����d�=dZv=��=)Q�>�h��8Z;� q:ǎ`�v	����>$�ܼ"N��p�V}�<hl���3=K(�=ؽ�� 8���P �Bs�=��;��M��Xό;�R۽奁��y���>=��޳�=f���H@�2LO=pi�=�{�=�d潵p���<�0nk�\'Ҽ��H�a���vH��*ս򈽈� �ZҐ����=��!=J�:=��Y�ai��,z�= ��������\�,=��=��x�
�yMB�x��;7 j�
z�=�n�=וֽ@�=��<<�_�=��3����=�IS��&5���=%o��z@3,̿6A���g�<�=r1��:��������`.>Ǎw��g���\3=+3��%!e�/p�>	0�Ǎ�>�
*@���?��=j���	��Q�����xr`�p�!�O�>��Α���=��!�\H>���=�vI?.��>r8�=]�">+Z>ͼ�$�=��G?B�c���V�!2T?L�>��ս�#Ŀq�L?8��?Q!,�a�D����U]�<λ=c��?Į�� ����ٿ�y=�6�|?�v��8@�NQ���T׾z�>���>�O?�8�=XD�����7�~?�L����?ѽH����e��BC��]V�?��>�@��O�W��;J9@@>��X��?o�$T�磿?%�<�r1�J�T?��=��3�Q�;����=�m�>�%�0��=}DC��8.��Q�(!�>�?���='	�?yI��O�c���W=�=�PX�;懙?+>��|�T�:����<40B�ז!���@h�>�*���	�=h=���l�(>�O�?.7���� ��N¼?�軠�<T,=!ĿG�Ҿ`�����>/=��\=�X=�W?��~�����?}�>��t��~��->�
Ľ��?@�d=���� ?���>K��Z����Y	�v�߽y��0����U�=�(��	c�0�9<d���� �c�¿�Ⱦ�nȾ�7r�jk�?��8wt?2Ƚ��t?��>A�6��U7���>��H����=2=M�V�I;���G��4���\�<J���؊�0��<p%��C�'�)��>�r[�0GҼv���,�>�jξř>>s�t>�y�>��Ľ ��R���=W��Oֽ%��>傾���>��i�%>Sa����_>��P��9�F0J<Zk�>o#�ظӾ�,������9�=H���w�ܼE=��=��&:�>؝��|����$Ӽ�xٽ���>���=�=�%K=*�>u<�>$���wu��;��,�����p�X�kZѽ��>k��;�~v�ؤӼT�=��s�����O?���uFe=�����[?�-�������x��=�r�?�ž`��?q��<����
&-�������=�ὃ��p�>�a?����1��Í=͹E���!=ˆ>p��>'顽����]b���<��5��/�����=�=X5=|�Z��K�="k?~H*�m&��-���A;>NO���)>^4����=<d�kDI���>��ܿ��1��N�>��ٽ�����m��̱?-�3��,x����=�A0=AmZ=D/�$c?��|�n-�`
��쾽��B��pϽ�'¿�쮿��ܓ׾9��N��оF�<���aO9��gA>�Ú��K���� ��%�<�;�<��'>���>��?1����3�OG��O@�Mj��Ž*�e������+	��o�>Ŕ5���\�6U���LM?�[6?^�[�\�E@��O��6��&�>�g�?��=kR���~Z?`$/���!��9�+��L�l��J�=��G�����:dH=|�
=(`$='m��r��گ�9Rx>�}����[�aJ���<	J�1}�3D��զ>!q{>H��>��F!�K�����`�T�j�	�����@�j����>:m�I�b�KO�>R|9��#>��g?����U�k�P�	�������AF��*���'��ܞ�:#�=�<?���#>�ߓ�A\�*">��^�a�<�=zK��f��>�Z�����/>��^@3�G𰽂I�>݅�?A��=6��=*.�u �<{}�|D5?#֙<��M�(�4�Y��B6��y��&��:!=��ڽe-ս<�=�p+�Su=�]�<(Q����<<�)��Q=#���L ����<�C�����̜�=佗<[�Q=J�Ƚ�&�8��&]-����=�ʻ��6���H���2�|��=8�<�4�=8��� �;�Er<=".=��}��`r<eg�����׽Lτ�/�ۼ�/��H��9k�4�g��󮽄� ���X�Y�
{�=��3<#c:=S��B� =���.ݐ�ĽĜ���m=6&���V�;f/�i �>��=% =O���o��N#<�=~�\�c(�^���Z����g=��l<���##�=��S�poi��D�; ��<X��=��\�qG\���C���R<Zy(<R����ƽ�K��iV<H�O=��<P�h�34�a<b����=�HV�}���<r$�=g>(�+�ٽ02��N�b��ټ<����=d����o��X��M%��Nw�p�$���~�Z�߽GNӽ�$��$2?L��?�4?v�Q��c$>�+̽�f)��N?Ӧ�>���?�N?�՞��;���C�ׂ�>O�y?w8�J�=��? x�>6��7cK>7<r>�"?�0&@?�(>M��?�A�?�}��*��>�Z��b�'��^��P'����
�?L?gȍ=���Z6@�*?�䮾���=��w���?� �?P��_��=��о���>S� ?Y+��p8@?
�>���ý�3���龠�?��������� ��¾��E�>�d�cg�>i�V�m�>�G>�]t���=<����e�_%.�񅄾ע9>E�?2�=����1���9�5�̼w�E��)n�h�����>����n>pF:�B4Q�ާ�;g�>2��r����ؿ�6���Ľy�e�&�c�]n�����<�1r=��8��+�=0j�>"�P<�jo�I/z����=�U>󘚼DЁ=N��=�>Nx=*"ý�񓿀��B������0��H	>A��>^��=^�e=xS�@�｡�=d�V>���>#ۦ�LYM����>$�=lD�=��x�}捿Կ��������==���>|�WP���=��%������e��dĽrL�/y?!G��C�S>;v8�Tٮ>5T缉��[�]��߭>����=����̻�� ��n��=�T5=�q!�|��=�T�����>yۺ�F�<��ýƐ��1F�>��Ѿ`��~߹<6�+>��p>�sZ=;��WJ�>��N���=����O�>l�>X\��v�;��ѽB �=%�}��'�>}=���(����(:d�=\&�=y*�0�=x�[=f1뽾J-�L�#���$���Ͻ������:0�������(��Z��ۍ������=�k����W<��=K������ɦ'=f�=�k:v�۽�H�=���Uw�=�M���o�=c�v�<Hw<�Q�É����C� &��y3	�S<�=����#K��<�<��;4�������]��m�=�U�=�ֻL���.BC���;D�>=�+$<#_9���ս8!�:��%���M�㽵��=%�����a�<�ǿ��<&w��YE�?@�6��:c�6��x$��zz>��Ž��'��h�����?<�M?>'>>��>&��Mq.=�`�⾧駾��"��wF?��F= ��0�d�z�t��5����N���L'_=v��=��}�����FC�wQF?�4p?�����	��Fi�2���`.?f�?�Z��(�\?k%G��T�=���=��y?��@Βn>��?��= 1d=@����V�B\ ?�N�<�����-V=���0�� �⻋�Խӳ��O<#XA����<o&�������c��-�=T�ɽ�oŽ�Q%=�]�<F���i�<�����"Խ�z�5B��]@�|м9����wϮ;(5��n�=!�ݽ��ӽ<�='(�(}�<�bʽ���I�����)�kSt�!҂�Հ�<�����B|��,�t*m=~X>+<���.��v�1�8=ut�p��<���=St7�/�>{q�0�q�8Ey��3�=֫��d總����v���~x��g&���"R>׼>�
N��"�Z$?�]�?�;��AH?_�_�.�>�&P����U=6����>���c���W@��A�ۋs>�i'>�!?��Y�3��>��k�^�?nO��;��0��<��x�O�~� F�<r� ?�"ؼ�K����)��pO�}��\G��K�;?w��> ��=�0q�n���%[�b��+߾q<��jc�f�u��틿��E��q�=}x�?��?���>zqZ�:$ݽ��p����?&=�>�_�?S��2�ڿM����?��ˠ�(����6�U�
b�����KU ?�-���+��>�X��g=����\��dW^?<�0?7��>����>�@~?�r*��4�=�P��mt�p�^=�q������,9�)}d�B����a�=����L���������>w�/?���؎>B
?e뗿0�B=ߍ߽1�����0?	L�>ym��ve?�8*>�?������A�+\�>Y U<:F/� 6b<^��=�� ?q���,I?=w�06�>��;��D?�Ey>}��=jK�텨>u��?�Z��7��?��ɾ��ؿz���m3�0n�?�9,?�*����A�?	@��L=}��=1I?G/�{ÿu8�W�=�Ic�ax�=̖�=4��)����=~�>9������˵A���"ڎ����>՝q?Mt�C�?�����$��ӽ��"$?�4p?^�=��S?v9����z���?�@��m?�:?P�(<P���~n>^�����m?I�X����Cg>=�ܾ^ap=�%Y�.ƾ��������O�>o1|>�X~��,��}��!d�J^��Xl���6��pN���>Z_���e�>��/���=��=e���ν}Џ>#�~���<�ѽ7��CP�>3����[�� �K�n���$\�=?W>�E����b�E��p��4�>�����νp�A<dý>�{�>�?m���d�<���I���=�_��:ͼ?����>Pa�������!
��N(��-�wz���	?aQ㿫����7?����6=�U=<z���$~�#��=�&@?M�L�ч������2f���ѾdS>�B>ʜ>���>�c5>�r?�`D��>�O���������#uN>�Ѿ߈����=���`����κ��>ͩq=�Pn<�cJ�>"��Zlw�&9>#b۽&������>� >i�½ �ʼ�A>��=���?�)F�$���[W>���=�s=�N5�>�,��c>�Hk����8+j����&��=��o>�U��:���kvz?�x�>�%��TL;+�?�[:�?H̍?���? ,n?�
���60�>�)?�-�<���=?��5�>���?�L�F���!`B���:��C���?x�(�HY�>_#N����zU=�1;�r���6�U=�G�X#h=�v���T����?�&>�����t����=��cTM�Ju=�.�=���_k��9>�!����=�{��>�?�=�埽)�>=��?U^�f)����=��=���F���)��?�پ��=�(�
T�>�Q?�fĽ����躒?�����?
��$�׾wil�J���Ƚ�>���Ʀ�9��?j�?�<+>��Ľ�}?�����G�#h�����ػ������Θ<��4�]�\�kyD=���������>�%��~XO>�.���i;>r���]��ՙ�� ������>����g>���>󫛾s?"1�a3A=��M�N�?��$@�P�>���=đ�=��s��=����N�?h�(�U� �I,��]�9?�;�?��;VZv���>f}�?��ھ�݂?��|T����>n����_�����ҿ����U�?��F?�D�=��������B?%����W<��a>i2��t�>t�6=������-���=�GV�����T~�=��<�od�=w;��g�<�<�>k>9#�>�|������W�G����K�>>G$?F �N�K=����_�D��=-�?E�?��C?�~�>8yܼ���=����j1�6�~?˸��Hv�>t��>��
?F�=;@�����6�>��?�J�?�?�>�A�����澠tl�;�N�C<W��l�>T %?��>�}�=�J��mp='�>��
����=q��<��.����<x0����/���)�1쐽�=�=e}�<� 漒��c�>���$�]=�e��_�
���>�g���*�����<���*�>��;|���l,�������=h
>kJ`>���?���>�L����=�]k=Z\�r`R��Z~?�8��꿽ͿS>�kN���=	�<��L��m����>%� ?k]>���}��g��-�K�a����@Ԉ�]g�"�X?o�=e�1>�9�j��=Φl={\&������?�����X0=�۾+T�w:��\�(�p�<<��#�T͇��q>���R���i�m�7m%�s�>��<�oѽ�D&��F%?	��>�ij��0&���5G�0���h;��a1>�C?������;銽8"�=h�=-�=��?f4���u�lE>�??���>�o=��?� �>j�>4F�?���o��[�b���Ͽx���R>㤿�*=�R�>�F>>j����=��!��
A?Z�I�*�hX8>�	Z?��@�	�<�@�ͼ	�����>���=�����=���=�5T��vC���Q>:��>$/ھ�Sj>ͥ���G���4=6!���O���V1>�.��P�>>蕿�ob�;�
�<J����?I>�%r?�����=�������>���?�	R�@�T@�����8�9�P�O�k�BԸ=%�ʻ+��ID�>#��>�Š���4?T���i�>� �=J#�� ��J��?���N�=h�>ZB�>�?��8?@��=W��=/n��⾞�B̽�������Qü��|���_>�X�����<o4?x���пlF3=����,�>	���V�~�~��='V����y��i�>�8/>ܕ�?���>Ha�����=��@����w:��)3<?� �=D
�l�2@YQ}��z�>a����0��zv=�78>�Ϳ�[�=�PD�������XH���MG�R��]���_)�eܕ����]��6?��Ͽtf?��>��K>>�.�B�F?m9�=��߳=��?�E�9��c�:(�������G�=���� �I�܀��Nƽex�=�8�><;?��=��J;�<���׾ |�<Si`=V�̽��>�$�>��ҿw�L��sڽ�����û+��=+�?�K����.=�,���<�2G�_�J��Hc?��2�κ��� =�����N<6Z�L���)=��n=C5���Tp��N!�(p��pܣ�+c��q����4I�������(�i�X��0�Xת=���=e����<'X��Xջ�ҼI�Ӽ1Ds���=jD��dB½�܁=����eL=8��=(�8�W���\�P8��r<�˼`�����= �]<�o ��[�4�齡��3���o����(<�CὨ ^���=.���鶗=X&�<�͚<���>�n�(^u=�㬿$�>g�?�!�=�N�>,�弅����Ѭ�i�b?%� ��Ҽ>����:�,���'��">�{=��>!Z��M>i��������>)�	>!&��
k�(���j~�>}2��>��:U=a������	���zI=G��=�#�=t39=�!>�kZ�����s
���pG>�?*���\�I2Z���?�-?r,��쉿?�Y��>,Br<m�)�%i����>��l?"r�=��=��l<�����2�?+Ͻ|������X�\;���/`=9ѽ���<�=<�$����=���*�̽�ƽ��=,�4��A�Rޒ=�xԼx���ѽ<G��]�)<VC=n�^��Y�<�_�=O�?����<���=$Ո�Z��=45��������=lW���q9��]=)b���K���Ƚ��໠�=�K%=�s�<�ݼ�s���=j⎽[���(�x ���=<��̵~�SE��_(k=�7�=pԔ<�2��t�@���N�(�,ӿ��>(�<o5�?@eO;��>�yӾ��=07ҿNʽ�f��po����B�;��|t�?��O?��Y>���@�����E�Y�0�>" >�擿��u?6f9>p�y�DV�;>L?ؙ�=`�r��� �[>L�>�P�ڋ�=�E�<r$�>���/ľ�3p��w¿BE�>����R����=Y��=t��2������JI_�O��x�W��*�<S���E⾜|��YT�8�K����="m��Ea�.�=.���92��?�=�m���D^� 9K��������/�S���{=�E��h�#:���|ŽB'����k�����ڽ������H�SA9=�SؽDn��F׽-a˽yR<����&�Ƽ�^ڼn������i`�Л��RA	��%=�T]����=����A��<�g����<����⎼�.�<�v���Ņ�U�;���P�7�7�{?��9r��-����(�;&)�=K��o�\=��=Tu��"ݢ=V@��;�=����TA�;��=[՘?@�?��E?�H�>=��<�{#�M"?��?^;��o�? ��irX�b���˳�z�>�-����	�ۢH?1[սT�?o�9>"�����>L�ҿ�[}�BӖ���>V�����Ͻ*{�=7�E����>�=�,�+ ����N=�qg �dv�= �辥�?uYv�o[k���	���<N:��F[ʿ�ڝ�7p�>,������D �6�=�$�p̛>�ϰ?��?�1> 都���=�o��V���s?�8�="ʽ��_�x\�>��=�?�<�`ѽ��
=�{�=�����F�=�Ge���<���=T�=��̽���nؘ�>���D��=Z'����ȳ�<�5���=���<��	+y=2V��8��|�ƽ���=@1 ��	�������~r��F�=8��M̽4��hX����Ƽ�ɺ�ߔ�=�X-=��I��=��j=ԙl=)�*=�=o�ҽ�C��^��$l<���=����R~�n.��诽��!=��=�*>��˽b ǽ�W?�	�Hɵ�%$��6j=HT���َ�$����#�<Ygl���m��XW=��������6?�d�˾�@R�ܽK�[�:�{�j�<��u=�x������+�"�b</j�2���-�=Q����+�<vX������=>�f?0?��\=�IǼn7��)������?�v�>�zͽ8�\=���D�?��uL�=���&�A��OG�?B����0�t�{�/Y��\�=��m<������'=읪=�^%>u񉿕�3=)z|�>���f(�?��)?.Ъ?��H�����X>���?7�>��?J��$z�H�8�YlZ���>Q��<�q@>����C?8�>w�W�ZIh?0�?(��>�h[�;��>lZ��l��R�`<M���Ҿ�=C��%x���C=�Wl=���=C����<�>'{�>��?>L����ѐ!=���KB?^r�=�~ܿ��M>rP=~qK�1� �Y���I�֕=E�>�O�?]z`?������xT鼈v���=w>�Ou?���?\}>� ����?�Ph?)���j�8��>�?*��=�?ҕ�b��JF�>*�I�ڒ�?_�>�J辆���m>-�0@��Z=��*=��}?Ydp���;>ϭ��\"�5����=�<�_s俴aU�M냽3�2>�EþL>�}¼T.��	��lɎ�=@T�x�Q3�>����\A?9���=����A>�U?}-�Q!��F��d\�E�h�B��~@��.?0$�?d@��L������x_�s�R?����Y@B"�?�N�>s�����<�W����=ʒ?�T�?���>.��=��<xߦ�-Y����)?3�C>���x��=6¿=;?\��>�S�|ٞ?�����>k�1?V�?M�v������<�"Ѿ��yl�f��>�����e�إ�==��Z�￀���\-�H$?S �>2@��j�?�ƽBĿǖB?������;�ѿt]��nu�=nb��jS����>I�?ק(?x��<�b��yE�F�8���?M�>$ྠ&8>X>��?�S=
�����7��>֊����?1��i�'�/8�i�@.��?��>JW�(�#2H?d�>��;�_�t׌?��?qJ7?$��>BF�?t+��)_��ؽC�ͿQ�}�$=��<����d�<�>�=^��?D�n?�k���O4>�֤<;�?ޞp?D�f������Xƿy͒���f����֗)�I�"���� ��=�]@"h�?�1��߾�=8�ʼ$��=r��>S���#�h?3�ν���PQ�����Z��<�=\݌�0��� �8⽠�)������Һ�F�
������H��<@����w�
�=R�����𽃡����<^z�������=���;�>=��w�d-�����(��=v|�=<����o=�C�� v<����n�&��H�����(�f��M� =��(�4������{�ֽ�%�N�����<`���z/�=L�׽���d�����!���<b��=��M�Nͽ�H=�M<
F�>o9G?ox�>!*��΋��{�=Ϳ���� ��>G�?�U?�����v�z����b>Ԙ�>�	=��0>�X��<�?<Ox�%�=��i�>O�?˾+�佬Z?˾'�������t󨽰
[�<�v? 1t���}��U��<��8��R�==��_����>����<=A9ۿ�⽪��=�AZ��oþ�%��B���K�:	6?ǝ��p�n��������S�?Ǒ�>�B����];g�	>�����o6����I�=a?w�����z<�?,=o��t'L��?��?B���[?]~+�lĔ�#��5�{��Y���f=)E�g��=����B>�U��F�'<QE>�uݾc����B�r=*�q������zq��DB>L�$��i<ܞ����=��u�6��Lk���?m�>��cII��}�<�9=�D=���>�C�!I��x�?�U�����<��T=���=6^�<�l9?bH��V����<(����/f�'��B���у�1\(�B�>�=�����3ǿݯd� BI<�Q콰0H<������P=�r��ii?W",�ӣ<���Qё>��	�;�[��&��٥��8�M�ʽ���<�]ͽ��>���σ�>���
�|������{Z=�׀=�ޛ�Z?=�v�=��ԽX4��&�?�XR��5�,g���T˾±D�j��=�o=KR��6�A<��4����t��7����=S��<���=pнbCӾ��=>L��s1��cp�5i�=�b���T����>�,?�` >^�<�+��K��!��?�$]�8�?c.��	;��7?v�w�	<���
#>���?�[A?���=��B=���A}>S�Ŀv9�+�M�=c�����}�<��;��`�ۛ��hn�W|����$w���<����?B�,>X�P���L�v��h��⳺�&4?���g�ӾO�u���>l?��>[����J+������AN?��?�y�>4~�>�J/@�h>=�u�x�q?��?�3�>6凾Nܽ��#�=��1<3�c�Q�n�hE���B>��l?���9Dο�wJ=-�?'�U�G�?�>��퓿��a?C����=x��X�; �FU�>�q;��d?Z�`�E�~��n��ԛ�Ԫ��@w�=4��M�=�[�=��I=Jjh?�u@>H4��>�����`F�-�=���Mt�=YH���<x�m�� ��m��0�=���:Z���9�>ƴ`?�4���T�=�Θ�L�5=i�E>�,<6Y�?���Қ�?�!�>�e�>v�#���C=������>��l?�z?�*�>A������!��3}�����>�۾�Kؿ�m���t�P'�?xXn>�Vg>RBc?j%��V�=�ˁ>��E?��0PŽj�=I���P�
��㓼�/�F�-��=C1;�R����nO>:��)}a?G��>	ez?; ����=�38=��@��y�> ��>����U^?@ꢿ��R=ӕ�=>�>�;�?�]����>�l��(@�=`2��i8��.�?pZ �_"*?�UN?�8<?Fc ?*X�=NĒ����=!�?%����_?� �N/�&��(��p�? ?�����Æ?�s���=����zf2=ˁ�>'庿a�;>�ǿ3g�>�򞿰�,?�M�"�%����0��=�,�>Z���P9>���"A��͸=�@�:
=��,?zp?&U�v��ȹPb����G���?��Q�� r�8���&`�<�#>����\9@� ?��Կ��b��=*�_��z���m�?Э6<䘩����=�VC=�z:=�5W��"��(&��<^=����v������r�1���PH<i7r��ߦ��=��<@�;��d�n��Ԥ�F"z=@"==�9[�(����t�<~釽�-��0w���y��3=�;�xO�xߙ=E��0= �f��Q��q�< q����=vB�6��=�[�� ��=�|����;�A~���C�7!��WЙ=�h���W�;4�=����Z½8��3���d=��������Z޽�O����=�(���TؼXm�=f����罿t�-wν�����+���	/= ו��&�=@��>%�񴨽o�,<�V�<~�-=���=�Ľ�U�������=�h�� ��<f:S��l�=|�ҽ0�����~�C{��4�P1�=�E���<�=�ȅ�<x�=���<G��=ܰ�<�'��!�=|��� ���h��<?=L)��⌷={`�� Fݺ�ys����= 3��$U�d��=S�`=���2<����:<r���ԽK�����<���͜�=(����<$1���rw�q�<�B����J=���<��A������6��=��˽D�<=���S��=���=K�b=G���H��+,[��M���<6�s=n����e�x�=<(��`�< ��:��"H��ȟ�= 9�=��׽�R,���㽱'�=ƣ���ܽ ���,�ʽ> ���}�㬽L,�;�k��L�O�?��=��s�0�T��=���\��ٲ�=��K��=���Cj��f�:e������<}�����<��=�s����l=#i����+��~��!=¨�s�=����O��V�=3>=�f�����=s�*�"���<\����Ϟ��f<�(<S��.���α�=�T=h}�����@�7�е�</�F�,��=��D<���=9��=+�a<�~��ܦ�����5I�<c<���t����k*%�Y�Ҽ!1���6��&F�̂��l�H=�d޽{Y�=G��<)����=>�=Ի������<�s
?⋛?ʽ?��_�e����=����^��x'^?�4Ⱦ�d�?��'@t��� ��?<�x��6�>�)�>3�;�<�<�	\L?4�Ͼ4�=g$?��Ѱ׾�9�&�?�%���"�|���4֖�[��7 @�����7>J]�ଝ��w��
 ?C�>3ھ�b1?�?K�W??L�ǌ)��(�=JR��OT`��{ھ�d��A�G>�3�>�e<{��O�=(>P�%>�'|��ٞ���k=d��?�+^���?�������i����<�"�<rҽ�.K����t��=�=0M���6D:�s`�=��<݀�<5��p�=S�"�P}I=wJ���+��闾��;�������\n����<C(�����<@Dd�3���Ǹ���=�Ƚt��=`�ż���f��Or,����>_?�n���U0���>�j����=t���c��l̯�2�S�_�X�þ�8��<p~m=��;��򽨁{<ܣJ��~h���3�ce6�{�%����=��������?�\?o��=�~~=-$��V���C-?װ�>�?25����?��Y�y�=�������w�G�E�T������?��,?��=�1�y�u�9��>��=Z�W>�B�PાJ t����c9ſ�v��Ô�=��>C�H=��<s׽c��>�g�>���>P���n��[��{?:ʞ;�Ƽv�?��}=3.?v燿}�)���T>�����=�ݾ��? {�?\�>@�p��z�=7�a�.c:>��\��4d?�X���
�?I�<���^-=�ʾ��M���<�Ñ�q#żvq�[�?���ռ���a{?�۽Ckֽ�}��ћo?�v=?,n4���!R(�N?����cJ�>�dٽ�r.���ｌ� =�S�� ?���=q��!Ҟ�,3=0���Hs5?pB�)hɿ���|�?��p�������=��t��>�<]ӂ>��=����Tt�~/?,؅=hK��V��>��=����?���<ho�<�*?
�����|���s�Pf$<U�Ͻ�Z�=h�۽h��<����_�= i�;�վ�dK� ��<�:#=V�l�{����{��B�O���"c��ޣ<�猽0hm=)GѼ"]�="b��d�<f����P�<��üj����,����p�=���v�8촽�o�<��(��{��r�i؉<C_�=��~=�x ��Y8���=���2=�=#�ܽ�=��9�q"��������6߽��	�\Pɽ^���:u=�d�`{��W�=���<@�w�$�*�?��=��?�˄>��>=$����ο�g��\Ba��I���2�(�{��UZ���i����=��⽱P�I@��i-,=��-?��Ͻ0'!>7������;؍�i-4>�Ĩ�z��>�%���㺾H޳<�Z{=D��K�=k
Q<pn���׽�ua��?���f�=��=O�%O=>a��h�i�h䜽�"?�C�=�0=�q�����\��5<��=S��:Y>RE���yd��e=�� ��=���>.P��9?�?�V���p�=Y.�={�-�8���8><�}?ZY��)��=颖���K�k���>\>:��>�[
�>i)?%���ƽh��=�@�B��>�0>5�>!����`c��m"=�⡿�Ė�1>����=$�h=Ьټt�=)�?�����mפ�%�_?��w?=ࢼ6l���!@�H��?�`i>YӚ>�(����K#�x��=���?�n�`W$>�!��'�=��=�9��V��>�ip�q>2V	>�P��E#?�$�>�� ?��=
 ������Fx}?�\V��E�?��L� ���x�
Y�G,<@��K@u�=��˜���>%@�p�=�䬿��:@'���T��?�(@��>X$���"@�2�ON�@G�q�$�=�7@Y18���<=$Nv�����Ț�m�@�Ӧ?A'��8�@f>�\v�����f>=��)V���p��i�?,�9����?~�ٽѢ^�3ҿÌ�@ng�>���r=,m�K�D����?�і?�"0���H�H3?k�>��>�������޸C���?��Z?�,�?�\s��д�Q2>0�T��>�/���L?'o?�">��=�����?�0�R��=f̍>_rG>��W�.A��t����Aѿ����^\=«¾ۙ��@;�=��U=9Ţ>�~��A���=dm�;�J���D��ӽ�&=i�A���6��n9>γ^�Vh�=���s�<��>uu?ZJ�?�M�>�i�=�	�=������L���?��D�d\\�i[���ƽ�D��/׽�o5��.���ë��Vǽ>&��\�4���=���<��K=�M����"����*=O :�߱<r�=L��d��=���V��Y׼4���6/�Ԁ�=�z�=�L��X!�=���*��<p`l�`$=@��=���=f� ;���H~!���ν �ƻ!^�� �a: xv�a���쟽E_��U|'�`����0[��H��n�=4���r���z=c�=Tfb=sG������������r?&C��b�>F��?ǽ����f��>}��?�Dv���?R7A�	vO���Z��=̿f�>j�{��E�;�ǿ��
@�&2?im�>�Qɽj1ؿ�rI?O�u1����>�j�R;~�ٽ���Ң����=��>I&?���=p���KR=�ٍ:4�����>�?�=:�X�˔ɾ"�J���5��z&4?�ap��*������z>u�O=Z��?�(@t��>WTc?�Q�v�ٽ��8l�M\�?����Ql>?}�?��/?�<����_���>�G�?��?���?�Hп��޾�,u���ҽ�Ӿ�ۂ��,?ǽ3?��M>��:=�2x�9��>L�r���+�;�� >?�=�j��d[=J-��`����;��];�����=�Hl�L�(?�#ʾ2��=�I�>,���c˾~ Ǿ���=�Ć=��w>�7B��,�f\���=��>���c�=�w���5 ?"
�?p��vW�=�µ��ʿ%���SJ?Ў��HI�??$�>�w"���?3��"߽�Ύ��gi��̽ߦ1��Uо�3�>�ƿ�̿��n>�{>>l�Nֿ%H�N�>=)�p㽙��\V���ۿ��軯�M�mX���f׿�X�=���M�> �ڻ�'�=K���_$���[�;T6��B��uą�5����?Ѣ�>�I?%�8�͎���]ѿ��>8>U?Ԥ��d���B�i�=���ۖ�^T��s=�T!��n�D����K޿�������W�?�a�D����"F=�՚=���vY�+V��h.<	��?��L=
4ӽ|��>Pni�?^ ��ǵ?x�8=���zLR�G���,�y�����=3�_��X><ر= �L�vT�=�Tw?������W=Vտd�=h�ʼ�&�>.x?���=U�t�W��R��t܋����>ɟ{��c�=U�>��d? Ƞ<���]�
����?���\�?�>��� �=,=pF~<���R�ӽ� �> �;�4�=ƧV��}�<,w�����?ż�ݾ2��>(�̵�`廈Z��z�?��=�a�>���7-��o���ܿ�|?%��ln�=Uϡ=v���bD?�(+��c=K�3��=��p?�?>}���[��<*D��%=?��=��g���>�J��ο��=ֿH�ۼ`���M?��C����Q�3?3z�?��e�� ������=���?���"���u*�{�>`���9=:��=���&6��fS���:?`�I�����k� 8�\�=^������A,��#=�;��񇲽�����῾���9?׃ѿ�v?������g�?�d=ߟ�<���=�7���9龳�>8���Z<D=����k��>�z?��\��Պ>��*��.ÿ ����j)��JͿ೩=�W>4�[���=tyz��ͽ���=T<��� ��?��?x���*މ=.��<BZ@�>�>��x>N�ſӈ׿�J�>+�콜�ł�>���>�f��p�оX�<�8=>�>���=?��>9��>f��� .h�H*%=r�Q�LBD=�"@>��L?'V�>�<�JZ<�D������`��A�g��s�>|bT�
X?�����3����Ծ*TԽJ�)?(�"��K)?�fH=(��>��=/�оTg���ak=��>˦��c�=P_��
ߐ=�) =V��=R�潷�6?TqͿ E��td���K>k!?���T������V���
9�����5��Ԃ��l��z�?�
�>��=�q?�!=�J������]��y=�<L���0Dd=�φ����=�ƕ���O��z��`&�^c���>�9�>ý&�p���<˦�?�Z�[׼3�v��ǈ=�i*�0��=�,�Iz�=M %���;����ֹ�=�� ��<دl=�{˼p,�=�"Y�X���x�⼰ة=�QY�I0U:�]=���+�ͽ��<�]L�{=��Hٻ�L�=���.����<ٝ=1��<��lP�=�Aۼ�G�<��3�E�	�'�:�����9�_�;����Cu?퍍:��0�hť�Qؽ,B���~����=��?�*�=S�?9�??�a�>ks>�|��=�����12�b���JE>�?>�8>�L�Ƈ�=��>%Ġ>BU@=���8��tq��@�c������(�f���)7�Lf�=:x�=b)>��p?G���l?��o�=�X�>~[R�_����=`=��̆7?@��(�=���D�>�eo>P����D���=�>�g�=]{�>.��=qC���O�˄�'�>3v���SU�gB��$Z�?��'?5V>|�޼��Y��>Lsr?l�ƿ��?_�>7@���?�|V=P<�?��)>�ؾ"-��u�@d�*>k�Ӽ���=mn���%@Z5>X�%?h�ž#�dB������!@�!�O��x>0�/?#оx�t��=��$>���G̾�F=�
w>��H�_����a�=��
��ƭ�h������?��k�,�i#�?�^���>�<�)v@��@�V�?�uX?���v��x}� :��4r?w��z뿑؉����ku�^����w�=`"�������\F�����MR�������G��`=~c��2�=�3w�`l�%?..��%��Y*>"?$�#���N?q��:��U� �4�4=���7�tV���%�P�ļ��m;՚��PI����>?Y]?��p���G�NvK?V ��j�h�ۼco���ֽ�b-���6����> R�"�=������>;�>ø>\�������=!�Z>��*����=a���d�-=���=�H�����<ؽ��7��F���~���*啽@,���S�<����IS�=۬��d6L=�P�����b��<k� ��;��U�J����y�h	Ҽ����HK�A�<�۽����!!���ƻ:6�=��{���=8���ż`�o<�s�=$8"=�^߽ =����=���X�����**=�Լ=r�d��\˽�=����%2=qĽ\-�6�i�X�xК=n��=���F�xە=�QM�(_m����>�|E>+ �}=����qԽf��֠���I�>b�?�/���J�νڐ<���T=�Ƽܾ�#>3??iBо �<�.<z`�=�;�%�K�lx:�ӂ>	���|�$�V=4d�w��Y>�v�<:򦽀�=�W<`��=E���1"�>�H��9���V�>W�Ӿ6A��`�=Ύ�=�nE>?���/2��(��>���/J��@�D=�~o�U�>���<�R�0�J<T�.�c��䂙�q[�>��>�(?r%�>y��>��?m�<�N"���?���?kh/?-i�?�\�/.�YK�����t�@�$?IJ�;=�m`�|;�?�8>h�_�h��=����޳���?�ڎ>�l%>Į���=E�@���{����=m�=���Խ���=}�=;���	�L?���>L�?V�G�>�% �g������3�����>US�?K����\���ݿn��=��<���1��?�٨>�i�?^��=��Ƽ��ҿ�W��/�?�O��/�NXt=k�н���< XM�`���鰍�ą9�Qֻ
���& =8G	�kT<Yk6=����6�<�z�<r|��ˏ=�����=�ὼ�)G�Xp#=�=�v��_)=?4�Q'E��ν�^�����;�����O���v���3<���3}�`�=b�����=B�#���=�N�;�=�%���l�=,t����ɽ�T������h񼨅�<����Ds=M�"<����:=𦡽2f����!�B�4�A]=j[D=d�'<ph=�e=�H�=�p��{��<��~�����U��,}�=�ּ�y'��F���I<����<��^����Y�<)�7���=b�	=~.�=Ug��U�н�Q ��W�it:��?|���Ƚ� ݽ(��<�1����,=���`�=�I�=�[����13M=w�:�O�Ž�@�;^�����=��'�u�=���<����!���#=���,ʽ�=j��O�� �6��G=41ٽ�OF=����c��ԃ= E�ƬP�K���>���/?��<�F��ey���̾~���|?P#���+�f�?������>�b����������@�� ?�^���
	� ��Q�?�y�s�=o��?|�&�&�<����i�+�>�2s�G;��뼖]�=z׽��Ms>��V?78�>��c?%����(m��2<�.&��U/�Ѝ=�r0�@��SJ��}#ῄ��=�ϩ�7"�?�:i?�9�H�+����<:��=����?Pȿ�R?��m�ǎ$���y<�VM>x!T=0C2=�� ������H>`m���м�R�<������_i.�J���u���G�=�;�z�9�E�'��ڽklܽ�^�����׭�I�O<RU��;���/����=�>������=���=h���4��=0��������Q��9�C(� ����������=�TY�2��ؔ�#��=�s�����=�!^��ý��="Q�(y5��s��u�,��K=6��=���!ݽ�@�k�O?<:=Q��?1I:?h�?	l���|���
����?a�b@�k�?�� �S�H������nQ@P�@p�*��-�=6�u�s%@��)>QJ+@Tv�?�����?^�@���>ݬR����4�#�����n��W����@��B���=i�F�����B�>�+g?7.�?���������<�Kי?���,����h��
�׿W][�O��x�C��0��nQ>�gt�I�R@�>/Q�?��콐&t<#B���3>Kߖ?��<<B����<$�<fL�Dv:=T	�O�=V�#���t������ӽ���<5�G<�J^�{7��=xt<<(��.�
����r�Խz���Ѳ�<Ed�ʓ�=/�E�5��Ҁ½�#սΖ�=���=¿˽����гR=�����"9=�̗��>��u��<��<?_v=M���́�tX�A�e<�J�<lf=>�u�nO�(ߎ���<���=,��OO���`��D%��?�=�坽���T�g�BE���#?���C����7=���>7�̽�_�M"�^c>2��?��q>N�	��y̽�H=���<x�f>�ſL��,d�?��#��^�>�n>�񵽺�d?l��>��ȽJ��?�����TC�=D���^��<��w=Q�2>`�N=X���R��=v�?y�{��E7�8R��8?
jo�v��b8����ν�J�/��>łU���俒{�B�{���C="��W+?��0?�t��s�>�S������.?m� �rc�>PK��0[ �   �  PK                      archive/data/3FB  Eu)��3��	����ܽ�C��|�;��>�����e�>�]��@�C�Z>�E�=Q�;_:?�i>/�i?b-�Z�?p�^����>����e�=���@*4v=G�3>�q�ϕ-���+>q��;�ƾH�=�Dk�ERν��!>��P>+�R����>"�P��oR>:����>��_=�~��*�h���?(	i���<;*��>��=Y/<D�d�d�<j�����p�b�?+"����,>Ay�>��]?��νM��)�9��E�>���>�q�>���\�m>�O����N>��<���c齴9�>��c��ߺ>Gi��!6�<���>kM?��+=� �/�2��h���c��(߽��*?<�'=r)�>�?~������>���L�u ��u�v�5�+>/R&���;��A_�/u6<?�s@��=;��e�i>�-'>��H�ڥ������o��~�9�׀���۽��D���Q��	$F!?�T����s�>�D2=��?�缦��=PKr��-      PK                      archive/data/4FB  ��T?���?���>�>�y6,=0�<�yS��1�<]�>~�R@F3<A_=�r���j���?jw\?�
Ⱦ��~<�2Ⱦ��~�����������>�M �F�8>+ �>ֵ�G�=S���l�?uu�?�p�꘢��|$��֋?�qb?2N��0_���7@�n<*7>?��H�?&P?�[z��m@��x@��?�z>��d?��?m�?s��������6��|?�>5�"��lT@��-��@�V	@)a�����=N����=�<y?!�4@��R�+\�t????���>7J<�|@�%��=�
m>���<a6?80�<S��?�W�?�g@~���K翻Ħ<yU? ��?M��?�"@)���P�Ѿ���@�4%=�H���N�;��=��w>� 
���j������ּŨ�>e~ƿ<�>��V��4A�i�?��P��ޙ��ݿf�?�2�q]�?k�=��>��S��/�=�Tz=(?�ᪿ�`������g�@F��" @�������85I�Ҟ?3{S�0o-=����X�M<�s3@�q˿a4����=;AM�VT�=���5@U,�?��y����=�=�?,�2��������a�@'&�>wm�=�h�>���;���?ގ?��@�,ҿ����g��ȫ�?�\��$��F޿�?h�ӺB��>��<2q�?}x�>����6B?pC@�_���<�'�=�>k@�P�?�3�=�K=�ӿ~�����>�M���W@�8w��?�@^~@Yg&��o�?�v��
M?Mo��ko?Y��=l�G?t��?��?�y=Z�'?�ɝ=�$?��<>��?��¼��b��p?���F����?O�=;GF�n=�>鉾2�>�2�?�׆?��t@�vw=���=BȀ���a�sV'�$|�<5���.�?�ơ���8�I I������1�>V9���ⅿ�����&�?��>/��[Vɿ/�!���I��)��sȿw�?�J�!v>�s����^� g����?�?̽'>�q��8�?�����v�=�"%9��U<�䎽<+οK��?�N�?�?� 9/=�g��U?��?%=+��)�?�%?LwQ�p|y>bo��G8=�O0?;@Յ-�y �>��2?���?zJ��-{<�q��Ģ޿|�JpL?�ڎ?�H�>�H?s�?0�@���>�'.=Ű�?�����~?�"?D�켼�׿���=�O����E>���> 
��ُ���ƺ��c��'ha>ў�>�]��|���=$ۈ������=�?Hl��t@��w?F�<+�?kG�>��?eiM?��>A9O?.�|�h��?�A<��?�Q���
Y�)�:��<@15@4�@?�? ��������ؿ�K����?�mt?��~��?�?����A;;�=W:�rU��gE�A�X��K?F�N��~�<nh?�C�?D�? �?��<�6?���?K��?�q�?<��1%P��!��}/�Bg���|3���<�_�>щ@`��xf����(���@��%@��=9s��u����k�Za�>�ܺS]D�8Gy�;��`Q@P?@�?�4l1=�� �e<
?tʙ?Zy��Rȁ?��?��<�x/�?P�4@�\�<lD�?L@ɴ�>�ڿ>�Qt����?X�L�4C)�w�>T�@��忐�-@�Ud?:;�H�?$�@�@��Ž��ػ9R?I�5�iS;?�M���s;Vd��6���v~��$?y�?E�����E��{��޼�:���S?2�;>L��{�6��ڽD(��cF?Z�����?>@ S�?���>�?t��?k�?�!@;~@�G�>7n7�_!@Ͳ��jjm@�m�9B߼?U�۽��� @<��?�@�@�+j@��<��?�&a�+	�>�w�\C/?�:�?�g	� P�������K���;P=Gs���g>�S�?��ɿ�~#��I >Ѽ�?:M�?y��>P(=�d��H��?Lt�>�^�Q�-��	@5E0?��e<�)�>f`��(����ֳ>��@3�<�9<��ҿ���=Hq@�Ɔ�;�\�PKZ���      PK                      archive/data/5FB  �G@�<@v{S@��B@PK�D��      PK                     3 archive/versionFB/ ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ3
PKўgU      PK          �od�p  p                   archive/data.pklPK          �O#�                   �  archive/data/0PK          ����                     archive/data/1PK          ��0[ �   �               P  archive/data/2PK          r��-                   ��  archive/data/3PK          Z���                   Ж  archive/data/4PK          �D��                   �  archive/data/5PK          ўgU                   `�  archive/versionPK,       -                       �      ҟ      PK    ��         PK      �  ҟ    