PK                      archive/data.pklFB ZZZZZZZZZZZZZZ�ccollections
OrderedDict
q )Rq(X   conv1.weightqctorch._utils
_rebuild_tensor_v2
q((X   storageqctorch
FloatStorage
qX   0qX   cpuqM $tqQK (K@KKKtq	(K�K	KKtq
�h )RqtqRqX
   conv1.biasqh((hhX   1qhK@tqQK K@�qK�q�h )RqtqRqX
   bn1.weightqh((hhX   2qhK@tqQK K@�qK�q�h )RqtqRqX   bn1.biasqh((hhX   3qhK@tq QK K@�q!K�q"�h )Rq#tq$Rq%X   bn1.running_meanq&h((hhX   4q'hK@tq(QK K@�q)K�q*�h )Rq+tq,Rq-X   bn1.running_varq.h((hhX   5q/hK@tq0QK K@�q1K�q2�h )Rq3tq4Rq5X   bn1.num_batches_trackedq6h((hctorch
LongStorage
q7X   6q8hKtq9QK ))�h )Rq:tq;Rq<X
   fc1.weightq=h((hhX   7q>hJ   tq?QK K�M �q@M K�qA�h )RqBtqCRqDX   fc1.biasqEh((hhX   8qFhK�tqGQK K��qHK�qI�h )RqJtqKRqLX
   out.weightqMh((hhX   9qNhM tqOQK KK��qPK�K�qQ�h )RqRtqSRqTX   out.biasqUh((hhX   10qVhKtqWQK K�qXK�qY�h )RqZtq[Rq\u}q]X	   _metadataq^h )Rq_(X    q`}qaX   versionqbKsX   conv1qc}qdhbKsX   bn1qe}qfhbKsX   fc1qg}qhhbKsX   outqi}qjhbKsusb.PK����    PK                     B archive/data/0FB> ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�#�?��i>0>�!�+��W��,�<?�`N��U?аԾC��?�*�=�m���:2��5����I?58��^?<#پO��?}0B>�vP��.�u����W?�ar�a�_?P,�W�?�i2>�o��4��0��&W?C
����u?�+ʾ+ʺ?ɭ�=0(��=��:��0�I?��'��Iv?�ע��4�?�,M>�9ٽ7[$�p?���%R?�_��K?䘾�~�?L��= �ʽə>������mC?
����|?����q��?��>>�ѼY^$�����T�S?8@���Y?���[��?h>�ս]U����~h9?�4��]?H��_��?{ &>ɤ</?(�j��
�U?u��GV?rל����?�RS>�!�����&���:Z?CD��<V?����8�?'�=g���y� ����|�3?uUʽ��f?��龿Q�?��>u�#�qF!������5?4�:�]?ҏ¾��?ɚ=���� 8��\����<?ޏL��_?^�۾���?�J>�4�y��⓿�!H?n�%��}?H���%��?��>>��/=��"�^Z����O?��D�73b?
����<m��>w%v��?F?�)���?���Û;?���zN==��>s����W?-d,��ɗ?ћ�G�:?�h���n_��m�>_���p@?Q�(��?��ݣN?qf��6�
=J9�>��q�<�D?�����?���3B\?Oҫ� ������>�Bw���T?��C,�?�@��\?������(=�,�>�Ƀ��ZB?Y'��Τ?aJ�Se]?cY���M�<Q	�>x؀��SJ?�!�E�?=�&���T?��¾G]�U~�>�{s��JH?{���+�?ׁ�)�@?����J������>?�{��fZ?Y �g��?|��E�M?����$-'��8�>�牿`�U?��3���?�K���I?���jH=���>%�y��%A?{'�k�?A���>?�r��ɼ<�T�>m�n��qO?�q���?�n���[?�[о̼7��>��x���7?��4�Qe�?���)=G?t��VY=_��>9r��qP?'z��Q�?�.����M?����	Ѓ=1b�>)v�x�A?M�'���?�!��T?b��R��;aF�>E$y���A?������?H&�%aE?5⎾�'>�ێ��=�y�>ϸҾ2�Q=����Ir������8>�ؚ��D>?�k�j7=�ƿ�W�f{���()>����Ǣ=^:�>��۾��=�ƿ}�`�`����k>	ܾ���=e)�>T��<B=Ϳ�mW����5>>-=ǾՖ�=��>p฾�0��S��Vg[�����.�='c�����<6n	?�;��q=��ʿ��r�*ж����=�M���p">NR�>�پ��=�[ɿ�L�X޷�k�>�þ�[�=a-�>���^��=�#¿_or�J8��->領��7<�n?x��C	���uſx#p�|ջ�K:\>qξ2�>>�
?Զ�ڃ�=�����N��K��ENK>����q	�<`S?j���<.����Bc����p��=W�ž�D�=�p�>yE޾ʂ�;l�Ϳo�s�tƿ}��=i������<���>�ؾS�׼Nο�_���¿�g>[���F�=�|?+��Θ=����?�f�X�ſhf�=IH׾/8�=,3�>Đ���Jl<��ƿ^�*���"Q�=���@��=j? xľ۽>,dȿ+�_��g����?ϮN���h?�� ����?�I?��=?p��?�t?���>��^�.rc?�}��h�?t�<?��V?��?�?��?��X��wy?Tr��:�?��9?A�G?�;�?��>B<�>��l�ԁo?,����?XS4?��;?�k�?L>?�# ?�T��z?��p�?�H9?!;?$|@T�?H�?p?U����?(���O�?~�6?��T?h#�??�2?c�K�;�d?��Ԯ�?��B?̻Z?���?s��>L�?-0b��h?b���*�? 4?'{S?��?�?��?wZR���?���׍�?N�B?�;?��?М?҅?iR��st?`���q�?��=?��H?6��?�
?0�?;0K�y�b?`��9�?�,?�X_?7��?�9?l!	?
-P�hq?�M���?nH??O0R?� @V�>\?�._���?�$��R�?$�$?F@?���?U>�>LT?)�P�tb?�'�.��?�8?�`?_�@`?�8�>|nh�A��?��?�?�&"?��:?m5@�.�>�v?��m���l?���f�?h	3?ҵ>?r��?�>�>o�>v��a��?��s�$Ȣ?��>������A�?	?�g>�3���Ԙ?�Mx��`�?h��>.��t�ʽ��?��D>�(��!��?Y�~�Z\�?��>�a~�j����&?��|>�ϻ�S�?�)r�x֩?��>s���ݲܽ��?@��>\��ED�?�S���խ?�|�>{q��h/#�]k?m!x>�9����?��y��M�?. �>2����o?��>�����ç?#�|����?���>-琾��B��?Q@>�����?�����r�?S.�>�s��Q�M�lx?ϥE>z�����?��t�T��?LN�>㪧��?���?���>�ۼ��ҟ?@���r��?��>[��������?͈>�0��M �?��u��[�?���>�R���� �%&?[s�>�8��皡?
z~��ߠ?���>M��1�X��%?�� >��7��?u(t�.*�?G�>�:���@�B�?��>l귿)Т?y�o�J«?��>��� ;��d?��>x���˦?+�z�X�?2:�>Ȅ�����kl#?c�c>h��cأ?=�n�$f�?̅�>��j��K�_�?�pO>H�?���?���>����-�?���h=d�S?��> ��?м�?�g?�A��?�K
��s)��a]?B[>���?Y_�?�A�>M颾�?G]	���=��R?��>���?���?3�?�瞾U�?�-�p��=�J?�x�>�s�?zi�?�-?b��h%?f��Y��.�J?,��>ԇ�?8r�?4�?�/���?��ޗ�=,t^?�gF>d;�?�(�?�o?�X��?y�r��=f�m?(U1>B��?>C�?�7�>����L?V) ��.=��^??)�>&��?��?t��>I2��H?Qz���>h�S?b�>���?~��?���>�Ͼ-�?l� �]��<Le?m4>\$�?��?�d�>�ӝ��d ?w���I�=&~l?�mI>B��?
G�?�	?��Ѿ! ?���)�=��J?VnP>^��?�H�?W?EQ��� ?�m��"&�=�J?ь�> ��?�H�?_�?,��?������<�[?F�>���?nL�?���>-�˾C�?¡�������Z?e��>���?:�?��>�ڀ�>����=(r?�F�sp���)_>U@�y�1>)ҝ�ք��W<�H�SX�ۈA�`��>ɹQ���>����ξ6�<�Vx��]7��eb�N �>%AU�C\>�U����P���Q���S��.��N�>�W\�$�}>_˕��	�p�>��N����3�𷅾��>�W���x>�᛿+��&���p���@���i���v>�U��8�>�����+��0�;�sDs�Ԣ9��o�
�>oE9�W�|>�4�����٣.�x�w��]>�A?��ל>�BY��20>s#��a���4�E�p�JC�h��Fc�>�=��,!>�������C;�Ww{���M�A9~���>�(;�l��>!R������2�1�p� �L��P��袔>�e_����>��徨4�a����F�`É��f�>/qO�~�>��f��jJ)��q���O?���
��>��U�i�1>�ܣ��޵@�f|��D�=Б�+Y>;<Z��eM>���������y*��s���N��|��q�>ٚM�'+H>�s���޾^>�/z��~iD�����q�K>��<���c>�)������2��^t�|n"�%va�'�{�8��=�t8?(�o�amn?��>���>�2:�7=�鏁���>J�5?�@y�_Yk?�E'>c�>��>���8���~��E�<0�0?��n�Ŭ_?��Q>{Y�>4)��e����l�=d�H?\{�-Nu?��]>���>�#���+�aሿ�
P��vC?�y�[�r?��>w��>�ˮ�q�e����?A=Z_A?��v���h?��C>���>�C�+��\z�����=��7?�+���MY?���=�7 ?@�[��C�*���&;��2J?�s��?Ri?���=�;�>�4��%T��T�������|:?"�j���w?m�=/�>c!ή�_�����\�h�p~8?mz��+wa?��=o�>؛)���o�(&{�6�=��C?	�r���v?��4>ٙ�>_�X�U�z�a4��΢�=~�X?�y�I~?U+U>���>k��3|�������=�!N?џ���$_?؄>y8�>91��	�X�Cᇿ���=0[K?�%q�ewf?��c>_��>4�P���C���z�	��=��D?�Tt�y
|?.'>�E�>�����4�?}���@>�M?�〿_�_?̇>	�>A/=6o�>�eÿ8׽}O���I�sd�?bT%�+/A�ub�=��k>�u��E�5��G뽂8�|�?D�%���<��$�=}W>�d��S���C� ��F��?�4�͌1��|S=�.>n�����������B.K��	�?���ױN��>��H>B�¿���~��ZO�H��?��9���D�>��>�̿�B�5Y�:bmM�,-�?�b6�K2��7�=��>vu��U���N�� f+�"�?,����:�G��=e�>>~/¿E$S��8�L6�+��?��7��W�W}�=��f>�廿ɍW��O��AS��m�?<�5�?�E���>�$>,5���S���<!+�L��?�m2�Ww8�<�>R�'>�<��Fg�b�ZY:��0�?�:�YZU���>���>Z�ƿy�Z��F��6i9�N�?@���TG���<��=�Iƿ����m���M�W�?^9���A��_�=�!�=T���K�,��_��-����?x:���I��d�=Vd>j����Pi����`r.�ź�?��5IO��6f=��}>�D�����X$�R:��r�?(����I��|��w��>�A�~��?x?��*+�1"K>��>�*=�J�����>�J���?0�6���ｨ�>?�>Q�0��?���g�>wP����?�=��qN�E~>���>��<a{����P>]wK��ݰ?2�;���u�O�~>��>B6�=/髿�V>�
<��B�?�h"���8�]d>�I�>`���󬷿��`>QVV�\g�?�U'�����R�>�1�>��*=i���P>�q4���?�m?�ן#�Ňp>/h�>�U�=[ȶ�1�}>��E��`�?���,X��(�><��>Ѥ=�i��-��>!�H���?���Z����v>���>���a���>i�P����?<T �^P��_�>��>L��o.��qY�>�&9� $�?0O/��r8��P�>4"�>)��Q٣�~�(>�)8�B�?:�=�$��� �>gD�>�F�������>ww8�P0�?~+��>E��>c>�i�>-���嵿��>�L� ��?�� ���L|>�h�>쟐=�,���E,>��8��Y�?4;@����pP�>�˙>UQ=�ߤ�Q��>��H�h3�?��?�ٶ1�Å�>&��>q��<�?.�P��P��<��>C����>�e�?�>�����
?n�Y�I9��2�>?����cv>EU�?g�>����?x#n��Ň��w�>�I��KIr>2ƻ?Ӫ�>O&e<�8?�fj�Ac���ݲ>�Ŀk�
>���?�}�>7�m��z?��h�kc���ۃ>�b��c�s>WB�?�d>ژ��X^?&Kl����4P�>u0ǿ��b>���?��>9E���?z8`��И�0��>u����T�>���?�
�>H �;4�?�!Z�7Z���U�>ÿ+�>���?2��>r!�<g��>�c��˕�W�>�q���!>���?�{�>x�U�P�?�0I��ו�0�>��ȿ?�>.��?��>V�ռ��?��X�����r��>3�ÿM�>��?֬|>�&R�B�?83\�#򖿠=�>�a��Z'K>X�?��>f��?��V�i�����>y����� >r��?;Y�>>�<f�?��_�Kq��|f�>�TĿ���=W�?8�c>�(
���?PV�������>S�Ŀ�cQ>�Ѹ?���>{W =�?�h�K������>%&���`�>Z��?���>Ir@��>%�ܟ=�zs���>{+�=�����>jڀ��>5��~C~=8ꅿ#~">�j�=r�����>G�����>#���\�=�ن���==���=����?)����>8�����=q�z�<��=P �͖?�����>�^վpUE>1k�Q�<*=^��/�?Ԯ~��z>�I	��0�=���ż1>�yJ=o��A�>9���U�7>����	 F=���_^>=>=�W�+��>h��)�>�$���>��q���<�V= y�`}?�;��AW^>���r>,k�5g�=��=Y ��>�덿4k�>����H�+>�y�+�=�B�=(�s7�>`��ŌL>*.�q8�=���o�=@}�=� ��?Xށ�S��>C�M="dj���=�4�=A��AJ�>�����U>���U7�=sd��>�^=Ɏ�=�c ��?����c�\>���6�W>���{~S=1S�<%��Q�?򝄿-�#>Sz��=`E���G>��=�o��.�>�}����>x��m.>sF}�u@.>,�b���!����>?��-�?�.~?F1?	kw>ؓ��1X�O=?{t�u>uk�?�U�?t@?+>~3�����I?��S��a�>w0�?���?�f#?�a)>85��AC�1�*?]Cr��g�>���?�r?�?�G�>����_X��%=?�~��	�>��?��h?>�/?{҂>�(���A�1�??w�G���f>	��?Ni?��-?�Vo>����$�'K?"�Ľ��>�϶?�vj?!= ?QRx>v7����&�I,O?Xf�r/�>�)�?b�?y�&?��9>, ��w6*�{�2?ԒD�:H�>�f�??Mt?B45?��>�����5��??������>��?��h?̩0?o�^>0k��K+ ���7?��
�-B�>�5�?�gk?��?y�W>�W�����Q�*?�u<��M�>?�?d${?�p?�uh>>k���� �O�;?33����>U�?sǁ?B4?T�>�E���O��UC?J���4k>�T�?'�k?�?Z�>nw�����L?�y��`�>o��?�{?�?Ga}>���3���PM?d=��H�>�Ԩ?�yn?�0(?��>ǈ�1��5�D?`�2�@W�>��#?k�?ᨕ?��?�g��.�?
T^��j�>o?��?a�?+�?=�>�ɋ�c�z?�t���?ё$?@5?kҡ?I=�?��?Y펿�qu?2�3����>�4&?�X*?q�?Y�?8�?K膿�v�?�����?o~?$�?��?�K�?�?#�����?����*�>#^?=�?E�?/��?A�?�����ȅ?O4��yB?K�?�K-?���?�v�?�J�>7����H?�~�����>��)?�0?���?m��?��>���u��?����(�?#?M?S��?�Q�?���>�ю�?�?sO��6��>j?��0?Yr�?���?ї!?[#��U�w?t����?/�!?�0?�l�?e�?�?~���Ύ?aϏ��O�>�=?�{?�ѝ?�?D�?�3��ac�?$�#�N�?j�?�f.?�u�?Q�?�� ?����?A����?t?7�?��?�L�?�;?/���~z?�_���.?}�?�?��?y��?g�?�x���U}?��W�j? �?��?�E�?�V�?o8?�HO�?�{x����>��?�'?T�C��:?��?֏���d?�k?D�
>�jO?z&?��2���9?!c?�����S?�΀?�>
�=?��??�R��C?Q0x?M��SO?�ۀ?���>Z�E?�<9?�E���?���?�u��Єv?<�g?�z>��8?�'?�%�|�;?Kp?W���*�c?$�s?ﱌ>�!K?p�"?_��R�=?�/�?ɇ��0N?0p?<wV>R�4?��?�Iv���D?bxq?�p����k?�W?qǆ>�	W?��0?�� �J�B?��w?%���|�V?J�[?E"�>C?h�&?x$���;?��t?�f��$�L?�Km?F��>��[?RN:?	�u��'?�tm?G����HM?尀?�z>{J5?�q6?`���n=?,�~?-<���_b?z�s?>A>RLV?
�3?��Z��5*?�2j?G^���Hl?�E{?��>�MD?��>?����!?��{?{��f�c?��~?;#>��M?�L+?��~�Lh1?��o?����Z?Kk?:��>�H?�?�OL���C?��g?����3_?z?Pr�>̃R?.�?q��
&"?��]?�'���h?~Vv?��0>�wL?�9?�SM>r��x�%�|�`�F�۾���>�X�>��O�2?��*>��N�<����P�����+?���>�1��E-?��>��H�����(�v
��&�?��?7�����:?Vq>�L�"��1=�� ��?w�>Bo�;S,?��=K��:�&���=4/����?;?"y�E?B?\"@>��-��b��WA����>�>���<?Y5�>��Nw ����r�¾>�?h��>���+%*?\�L>���!��7�<�����C	?��>�
�kg5?h�Z>1(�� �%����=0���>f��>Q���>?~�F>4v=��> ��E�=x�ﾧ��>	�
?lX�s�!?�~>0�%��#���7=�$���W�>���>���E'1?27>e.��v"����=���2�>[R?�%�"?��0>�e���E$���"<[��5��>x��>�n���'?d?>�O�� ���=�^����
?���>h� ���1?�3>�B�$!��W弧�߾=:�>��?�^��0"?�X>N4I��"!�^�r= �ľ�2�>˺�>u���Z$���@=v|�LM��>Nx�>|0��,:��t�>#��|�>�7�>�"�dG�>>3�>����*�<�ZZ�>�%����=�7��Z���>�Ԝ>����t��l�]>�#��n>.�ѽg*� u�>�>�沿v�?��Pj>o�"���>&Ҵ�����>6�>D;Ŀ��)��u�>3!�կ=�O��?O�k>
��������>��#�Ԉ,>J��;�p$�3��>�>.{¿��*� Ģ>/�VK�=�@:�_��� �>�P�>>ܷ�H�2��e�>uc#���=�OL��*����>hN�>�����>)�L�>� ��[�=v���hV��"�>ZH�>D�����8�*��>݅"�?�;=yﹼY��zY ?HG�>,¿��+��ϻ>a�!��[�<�(�b���>��> B��.�~�~>��!���=u(%�=���>0/�>t�¿����T>A���1=���[/�d��>�Ԭ>����F� ��mj>y�!��/�=ڳڽ��Z��>��>�2ſ���
?�>I3���>c嵽�g ��6�>*x�>�t��.0�DY�>���>� ���)�?�+�V �|?�?PF�=�jo?�1�?<u�>�V���#�?:QF�����?�{�=n/e?��?n�>Aݲ�;6�?4�Z��|	�ן? ӆ�؃z?���?�x ?�}��c��?*�8�l����?M� <�Qx?8ο?���>�}��7��?<T��p�d��?x�8=8�?B��?�W�>n���Mx�?đ/���pI�?�/�=v�b?�A�?MS�>������? XŽH���\��?�<>�m?^u�?!�>�g�����?3F.�l�ᾶ�?�M�:&��?�e�?��>�y���̎?J��� ��PA�?���<�cd?Ҟ�?��>Q������?HZ9�����?mCh=�w?.�?O��>Ὧ�O��?�g�N0ݾ"P�?��>2l?Zu�?أ?Eۮ�!	�?�7~���?�>�$}?"��?��?Ȩ����?����tN�P�?��Q=��|?P��?�5�>������?\@4��M���?��=�Yz?J��?���>�`���L�?�h-�2��趣?�~#>��|?�?���>�j���ތ?�:�2���$�?��n<z�~?��?�n��J�O?�¿�ν���<�x�_g�=�9�-�ȿ[����*?ۡ��(ぽ�O����#�þ�4ſ���nF3?-
ǿ���U�������>�s��k�տF����B-?!����8�.䯽�֍�L6�<��Ⱦ/KӿU���*?�VʿE?Ľ2�������{&=��⾦�ÿ�g��1,?9Ŀ�@��Žk���7�<����ARؿ𠏿��O??FͿ��-�NB�<i�s���l=���ɿ�O����<?o�ɿ�39���H��p���)�=���	�ӿ.≿by1?m�����"�Ԗ�7D��Xπ=tiž/�˿ ��� �9?��˿;3���_Խyi����=����O!̿�匿RBE?�¿7�6�7�/@��vi�=�f;!�οnm����??_�ƿ�����*�h���^��˾�JпP���.^6?� ��)Q?��
!���r����=fҾ�AϿn����|C?��ſP?��R������r+�=.Y;�տV9���P?��ȿ�	����<��y�k��<l����>ƿ�o��>�G?�ɿ��#�"� <�|����=T�پ�̿?����?Կ�=B���l�>����>ԗ��i��?;���Ǘ?�=J/���jG>˸ҽ��>@&����?�I��{(�?9��=Ř��U�>Pg,��>�>.���+�??�_�k��?�q>*1��i)�>�~,���>o׀�5C�?F��w�?qD�=�B�����>��+��~�>�
�����?[�p�qܘ?�>�z��7�v>)�ý}��>
Cv���?�Ը��Ϥ?�jg<����&\�>a��u��>�bn����?ނ���?w.1>DI��u�M>�$���>����b�?�k��k2�?�6>���x8>������>�?��]Y�?!������?UXO=.���Dخ>�����>����j�?㿊��H�?��>�h�����>�����>�5���M�?Q���E(�?�B$>\N��Z�H>浵�G �>�����p�?]r���Ǔ?�>����i>R����>,f�I��?�xV��?
T#>,����{�>�j����>P���s~�?�V���~�?��<Z���J>R��7�>���ǀ�?�釾�x�?�Ϥ=����M�:>��=�!��>��e��+�?�ɚ�o=���늿�N;?��>��"�D:�
��(��=�������׌��|$?�v�>�f&�� ��_ý-F>�A���{о�v��>@8?ټ>k,)� 5�!M�+xs>2硿�ͱ�f(��9?���>�,�/���½�,>�������?f��O�+?��>�����FK���=H8��w��e|���?蓖>�[)������ս`b�=^��|�̾���VD?���>-��0�!�Y۽uL^>ꛤ�<	��<���T=?lc�>m�&�2�:�b( �k�C>���t�������?�?�L�>�,����^�\	>�8��K�۾���6<?���>�m�`�!��aͽ�o|>�̙��/ž:����;?�I�>����/��QG��>*r��"���=��$�2?ψ�>m-���'��-��>EN���Ǡ��h����7?)��>�!�h��@4�����={���[;���,#?�G�>���8��_�e�/>n�g��!p��d�%?��>���>0�L'^���>�����z��Dɖ�&$?��>u����&��V_��<>��(�>'w���RL��Q)?����4>(��7�S�)�`��7�x>�ι������"?�ۋ���f#�-:�ǁڿ�D->Q�ܾ3�P�w%?�����U(��$��� �b�߿��?>���.����?ˤ����Gq��()����>;���~��Y�'?ɺ���G�9��Ϛ;��� ��>뱺�,֤�%�+?_����
�B&�:(��9㿴BL>)A⾼���5� ?1����{����1/���<?p>��о�S�(?������V���7<�ީ�*;.>!����R�]�?����+�"�W���d�	�ڿD7>-?�j��u�,?a���G%���;�.��i����>�w���79��!#?�;���:&��F!����IۿB>�>w��l3:�#�7?SK��+P��	��>��*��!2>!�Ͼ ~���?w�������	���A����h�>�9۾�����K?���1�����O>4�>$���
>!2���TO�g?-"������l��66��d�p9>�Y�<"�[+?O2��|�"���*���(��O??���冾)��W�8��(?؊@���>à�?8Ca?����R�Dj��Ҥ��?V|@�"�>�N�?��^?Q��������<�K,?��@�Ь>���?�X?*=��l�$�,��=��B�?���?n��>_��?.T_?!vm=4���<�EJ���-?@ɬ�>���?��[?�mŽמ_��C��C?��$?�|@�*�>���?��m?�Z�qpe�Bv�֐�<�+?�h@"#�>3<�?J�a?��b<��c-�������� ?ɖ@���>���?f�k?�&ýr1�?Ž��ɻb�?v@t��>���?pOr?Ukq=y!ݽYR{�rӽ�l?�:@���>��?&i?�_�<��O�d�&��惼��?���?f�>E��?��R?xBL�+� � X�������
?�@`��>2�?p*^?�'E<�=&��7<Q;�p�)?��@H�>�0�?:�T?j5N��-R������l*.??��?Vh�>9@�?$n?>==�=��c�����G��J?zP@4��>K��?Z%a?�=j<��q���P<���� �#?�& @r��>��?�x}����7;���>�<�^t���?\��>�C����x�?�d�;T0�X"�>�%�-~o�6�?���>�4�;R�e�+i�=!�(��w�>����~���?~X>b�����w��#�;�`C�HM�>����`�M�(?��Q>���<�{��J=�=D�� �>1)������y(?��>s�=�^����=k(C���>���|�{��+? �f>1�<"�U��7Ƽ�O2����>�Q�,�`�U,?�1> ��<̷a�j,̻��?��5�>�*��Kn��1?.sd>�����n����<�	=�tO�>�#!��k�׀'?�1�>�NW=�M}��_C=k9E�t��>;e���c��)?��>gX=R�v�Z�Ѽ�M�Fݮ>Au��ki�Ώ
?&9i>#ϲ�M*m�xY�;ѱM�4��>ɗ�pp��v)?�6�>��=�o�G8�=�G���>���ǀ�E�?D��>Y��<�g�4��=[g=��>U���t��?R}U>�\��` b�|>�=�3G�*��>_�!�Iv�n�	?���>"[����d���:=~N����>�1��cf���&?��5>�@�;C	�z��?�d?
�ؾK�>*>S=�6j��������?R��
��?B�?Ii���>�O���hu���>R\�?Ȫ��Z�?$�?+��K��>�C�2ku���>��?n|&��G�?J�?�
����>�s��-�o��<�=�)�?����	�?O�!?,�߾���>C><�Y��}�=��?xd"����?�?M�
�5f�>T�	���n�w�к���?`�'���?�]?Mp����>�	���V�|˃=6�?,�+�04�?2�?{�����>�q���Zq�T�>S��?.�1�`ٻ?��?�B�W'�>L=Mc����=���?�V��k�?�?!�����>��e�Z�Ƨ>EJ�?��1�� �?8_?��
�m��>0�;<p��|>M��?�v����?fD�>�־c�>���<uT_��� =Q��?&���t�?[*
?�L
�m9�>�C���lX�5d=N�?����Ļ?S]?O\	��r�>��_��]W����=

�?�V� ��?�y?)f���>��=q[g���=���?`&�`7�?��?�3�u?�>4���;]M��v>�C�?�Ⴟ-�q��hT��qþv�Ծ�@�?�b��R�?���!Gu��셾8�4���̾蕏����?v,m��?�����i�!�����U�U�ʾP֭�ß?{cy�O��?�F��&r�}����Z�����o��拫?5���_O�?���-��~끾l�8�����A��^:�?B�6�Oa�?����m�y�^�ܭ:� �����˫?"�X�{�?��MTf��f>�(P�yo��矾c��?�D���8�?8����x�0 ~�NB=�{��^�ξ�?J^l���?X��k�Z3b���A��E���ξ��?��Â�?�L�х~�_Rh�)lN�����F8��6�?������?���=c������A�FO�5�����?��)�e[�?�%�{���t��G��8޾l�����?:��4�?��o�k�f���q/W�}�˾�⡾��?����Yǧ?�W ���p�^Y� WK�?�پ�׾f��?��*�9/�?&���_b��؈�b�6��۾�鑾N�?X�����?������f�r2��e��t���1;�?bB��ţ?nv���?�JǾcs�J���Ӄ?:�>��>����>��?���g���	�bk�?�1�>�>����r�K=�,�?^Q⾫C����2�?<d�>2M�>���L��=���?����)�*i��6�?d�>�>����9�A�?}���)��P��S�?���>��>5������=�Z�?�i��O�)�ei
�T��?Z��>��>J�ݾ��<�ƍ?Q�پ��,����?�V�>p��><^	�/��=]�?6+����
�
�l�?��>���>Р��s>+�?Ѿo����	�n&�?���>���>����>
=�ч?o�۾�B����o�?�r�>���><:
��%>cѐ?��Ծ������&v�?�u�>R��>- 󾱗�=�׈?�1��������Fc�?�#�>���>���vc=�?ͣ¾=~	��a�@-�?:��>M�>-K�-x�=a��?�Z¾� 2��C�pߐ?���>��>���פ�=]Q�?C�ھ�8 �B�����?�خ>�H�>�/辳5�0��?畾�$�Tk��v�?3�>���>�i��>�"?]��xL?��l<d��?�ξz����T?����9?�K���$?fݽ���?K�ƾZa)�ޗu?ȯ��,?�4��A%?��B=�0�?�	�<E2�h�l?� ��a.?��ʾ�=)?��v=�O�?��:���K?t��n/7?����i�?�ާ�@��?&����9���q?6U���/?ʘ���?�m=��?F� �J�8�l�R?�'��?V���8�&?��p�8��?�2�/�xbn?A7�Qx?����?�s�l��?���t.�Pe?e�
��?𰚾H"?��N�?�˾�71�
4N?@w�#�"?���C�?�ٔ���?[�þ�D$�n}i?� ���?�T��!�?���:��?���>	���f?�V�Ǎ/?�"���?\ݗ��g�?�6���>�D�l?p�#u?L����w*?����P�?�b¾��:��"L?(�
�o�?~�Ҿ�"!?rȽy�??���,���Z?���?�g��	�?�Ͻ��?���8��\X?�*��!?������?#�=V��?l��$���\?��o�?nP�dd<��8Y?\壾d��>�C�?�H6?+�?k?Q=����QS?^���~0�>�$�?Y�2?$]?Gj�>�����G����7?/Z����>z�?��?��?m}	?�7i��A,���E?A�����>-�?�t<?]a?+h	?#�����<vXQ?�@��L��>��?��2?q
?�?��=ɥ�;��Z?�m��̆�>�Q�?cN3?�q,?@��>�ͼw�ݽAW?�����>(��?��'?��&?;c	?�>�<����d�V?hQ���-�>�s�?˘?�.?��>�$����0,8?�搾b��>QL�?c<?A�?�?��@��';��;?.����>"��?��2?�?�G�>��=6�����L?�ߺ���>LR�?��2?�?��?�	��[����^?�$���%�>�ޟ?�2?�Y?�;�>ń:&�Y��I?��W�}��>�I�?ŉ$?��?��	?���=�LJ���F?v��R��>���?�;??��>e��;�ż�_M?0���jĠ>�%�?5~/?$�	?�?��o=�q½�9?�����>��?�?%?!B,?������_�~`v�?B?�xj��оF�¿���<�n�����#����{
?L^|��̼�̿!s=����/*�A�?
�<+T?L�{�D-��6rο�4�=�������a��ڡ<��>
�l�F�־�CɿD=������"��KO���
?�`[��Ϣ��ɿCS=���I��4�ͬ��P� ?�T��^˾��οuL=	�%�q��[83���<oJ?@R�T�Ǿ��¿��=t��	���U.��{^��+?�1|��մ��!ӿ1�=�U%��P1��9�S�Q<�"�>� k�H�Ǿ�Ŀ�d�=��q!��Y��=�?ȇh���;�1Ϳ��=;\�;�������!�A��>F�e�༪��+ҿ���=�<��/����P�����>�r�Y���XMǿ��>Ց��1�,��.���k?tOZ���ؾ��ɿ<�f=����t�U+%�����Q�>�u����Vpп�.=w�����]�2���ս�e�>z?S�]���/Ͽ�0=y�%���#��+(�(�=��>P{�.�`[ӿM0=�S����� ��٧��S>p���>��J��V%��C��9�þ&�
�����L2->�&�� 'z>�~J�?h4�N����韾z���՟���>1z�<��I>�`��N:��Z��Eb��B��\�����5>5W��»�>�{Z��#��Q��Cޙ�(	��VD�M��=D�*�9�>~F�٥:�"i������h�E��v
t>�EX��q>u�A��q@�
W��G����_�mk��kߩ=]��=ٿR>E5_��C�����9����X��� �j>C�=*�o>ǁZ����@���ó��4�d�4����=5y��!<>JU�gH6�b$��������������h<>N�*=��>��V�Cn0��C����l�����Ix��<�==�$��0�>3:Z�����������
)���q�2}S>'�=K�e>'�^�I%A� ���Uf����+�����=_#�=��>IG��@�d����	��f�	��>��&��=��6�0�z>z=�):�M���蟾�����L���>�$a��Ǒ>�&c�-;�詨�{N����	�������=@6=�%->�$<��*��c�>�|���U�?+?�b@��??����e>��?�O�>�r�R��?�U?�m/�:? ?��"�s�	>���?�ɕ>z��2��?$��>�J�8)!?����.�>�h�?U�>����,��?�?��"��]?�0 �Xc>ĕ�?~T�>��: ��?b�?*\4�& ?���>x��?�"�>������?�[?,E��
?�M��+�>���?���>�u�PZ�?��?��3���?".��/��>�-�?��>0ˉ����?PD
?�5���%?�n��%>�5�?$��>%��Ї�?pp�>&.���?V���C>���?ʦ�>oH���+�?�?��8��s�>g�߫�>�]�?ݬ>��Lz�?83	?��K��Z?6��h,C>g�?�
�>5�+�r�?��?Xp(��?>���6>��?p�>����dL�?���>>�4�%}?������>l@�?�K�>h�O�Ds�?���>vr1�"K?DZ�@C9>^��?ޫ>��I��I�?��?��8�D$?�:���d>���?�`�>N��RX�? ��><�'�T�?����l>@R�?��þ��>���H����Ŀ�T?ۘ�>x�m?������Ѕ <=���󓾇�ʿ��?I�>H|?#Y��r�ѾE��:�b��þ)�����7?��>+zn?�<���^� �=KP��4������En+?�͌>�Dg?1���ᘾV��=�� T���1��ib.?{-�>�~r?�ߙ��D߾�=3��vɖ�G���80?�>7Zf?Ԉ��#価�;mu��h���7��)�?���>��{?�В�^5��J��=���D ¾S���?���>���?)o����վ%�>�-�v
��P��w-$?U��>���?�/���辱��=����؅��a��Sj?��>���?�Z���};�a>�Y��現�X���K?L*�>��y?�p��"�Ⱦ3kP;�+��Xƾ����E!?s�>l�}?��~��6d�=Q���~��5>���t?��>@l�?�i�����{ׇ;Ƀ��ֆ��U��/�?ϓ>Q�x?����xξ�A=�T�����7�w�2?�f�>��q?�l��J��nm�<��"���Fǿ��?q�>0ބ?����6���F����Wy�>؏��$"�@���d�̾�'G���}�A�;��﻿E�>��v�؅ݾ�]���颾q�$����(�\�����H�>j>�����ӂ��{���R8�l�����>��ú�3��>l�ľ�������R��oS-�����Yt]��(����>�;j�&��&n�=أ���4��"�Jb:��9���P�>8���U���Rj�������"��]��G*d�J��c�>�'��D����L��M*������^�|����q�>��ľ��߾���e����>���{�>�[�h���k�>���,���+n�L̴��D�~<��BWJ�*��@�>��ľ��ϾA^����ƾ�iE�b#}�/V�6f��a!�>�~�Hj��<�������sK��K���
F�x���� �>�T����6���bӾ�L:�����Ǯ^�PY��A�>�<����C��0Aʾ)iD�������S�<��
�>ܡ��0��|e��^����;�����T\�,������> g�������Y��)��?:7�~����Y��ܩ�;I�>�Ⱦ�鰾����E���t;�𡆿±q?�Ft>e����>Y7�������O�����>x���)�?˺>?`���t?g닾Lr��I����>�a��w��?vm>C��|,�>5��إ�y������>� ����o?�Q�>=r�����>�rվgT��B�m�>(������?�s�>�~��\��>A���dM��#���1I�>����l�?q>��C��>�宾u���pd�b�>�|�3�?�d>��`���>Ox���x��.��>1�}���z?W�A>�jX����>;9Ҿ౾t6���>h����,�?\>��{��N�>�s��(�Z����߇�>F���:�?�
Y>�]c���?�ɷ�g빾S� ��ҧ>n�u���?y�P>��Nj�>P���&���(��Ð�>�:���J�?�Y>�IP����>��׾⩦�O$��K�>�ׅ�A�?��0>�j]�al�>�����Ts������>Z|�X�?�-!>X��!�>�ǣ��ǅ�����~�>����ւ?e`>�߂��c?�@Ǿø�]����>̷{�"�}?_�U>��v����>1m���X��a����Q�>a�z?�~�;���s�?��??ᄿ��X?)zm�� <Ղm?��DY���ʳ?3?n��u�J?E��������#i?Ӥ�<B���x�?PX?������U?�5x�a�L��h�?fl�\Ǿ"��?�� ?��y���B? -��j�����?_NɼP���u�?�8?�Ix�C-R?��e�,�V�yw?�TK��������?��?�,���3D?��x��������?U������*�?0=?�ڂ��vd?O3��
=N�U�l?�A���$Ⱦ��?�?cu����G?8/��
RG��fa?������þ*I�?��?��z���Q?��f��[��1Gw?>9��(_��L�?��?Z�x�OGL?a7k�~�n��v?ߪ�;�4�����?S�?�)y�g�d?u�l�j�ݽ��n?~{��s�j��?��?zj���WO?�?���[н �?N	۽fyk��ɶ?�H?$����e?��{��)�A�\? :��$>��\%�?���>�0s��@?7�{�Q	���]?�i��*I��B��?%�? fn���Z?7���䴂���z?_1�6���Hۿ?��?�'{�՜I?sm��Z ������?P��� �]Dq�6l��#�6?C�>JZ���w��1i�>_�����n���ڮɾ�/?J��>�-�����*��>b2��H迵ⶾ 8���0?qy>������ɿW�?���\����J����%�?�>׋��ǿ�?��
�L����6�������$4?�nY>zX��i��?�o �A�ￔ[��i� ���+?wm>���g���K�?�&���󿴰e�J0����?�À>�������-�?�
�#���s��ھ��,?��t>�'���oÿ!� ?���]@����"�¾k?SZE>F6��I��K�?�S��+�md�\߾�.?�;�>r����ɿ��?���Ǫ����.���Q:1?��Q>U��8�Ŀ�S'?���Y�a�* �ې.?<tu>�M���¿s�?ز�����Y� ��'?�Qb>P���Z����?t��AG��࿾�?^.?�w�>jY}��<ſ!�?���N�^욾����)N;?S?J>�Ӏ�����9�?ӻ�';�R��� ����)?5R�>�����>bܾ���?�S���ֽ筤?[~����?T�?�k�>����&��?�W#�o��m��?ո��G�?�&�?�°>�վ>P�?XM��͆<��?����Wύ?���?z�>��ܾ ۾?x�!�� �� �?����[��?<D�?�"�>������?�l�(B3=ģ?�CĽ���?�τ?�0�>�.Ͼ��?>���^����?��s��v�?a��?���>M�־���?����`�iӜ?�;0��R�?J�?O�>;�վ���?�(�� {��X�?k�轵˒?�L�?�v�>*����@�?�B'�|�]�c0�?&�ǽ
��?F��?Ŭ�>�t��\�?����wp�1"�?MU�v��?舏?(;�>�Q��~�?]���=Q�?�:��g�?L�?�i�>�2��J��?I�������?v/޽>�?�)�?���>گ����?�Y� ���&�?6'����?"�}?���>N��d��?��"��V��ߊ�?�����?�z?g��>������?)a�j;��?��ٽ�ϙ?�ׄ?��>#!�����?�$�˳ʼ�Ԫ?�-�RȞ?�֐?p]�?�g�<u�X?\�,�)�,��A��?�X�>��"?L��?u?=9T?Q�ݾ��2����%%�?���>� ?���?���W�P?K��ָL��Ӵ���?6��>�%9?�+�?���S"N?�MѾ�.�>�׾�r�?���>^�2?���?|����G?���n�9�"�-��?�~?�Z>?��?~`�=�Pd?�����6� ¢���?���>f 7?P��?�f<�X?�g��H�E���¾ye�?И�>��8?@7�?H��+IN?��Ѿ\A@� �����?���>6C?���?�B�=s�M?����tF�no���߿?��>�5? *�?�*>��O?��¾�1�$t�;��?,* ?��4?��?�x�=��U?(����?Q�����SR�?�8�>tY?X��?� 2;u�h?�u��|�*�������?t�?�:?�y�?~�=]Y?�Q��~_9�f-Ծ���?��?X6?D�?��=9KG?�U�R�?�jq྽��?h��>­3?�,�?^��<ѳi?��;�~0�N�߾���?�]�>L�!?�E�?
,�=��i?����/�.������?"�>�W-?1Z�>Rz��x?P�>���=$rT>����>~���Q>*��$�n?�]>��z>��>^k
�S'�>mJ='i>�@�<�߀?w�Z>�}�=+>c�����>[ے=j*>R�����?�5>դl>U��>��0	?`�
>>c;>��t�{�?�n2>��r>r �>p�
���?��=�$2>La�<���?���=��v>z�;>����v�>��<��>� @�� o?��=�'>�u>Ǿ�<�?��={zU>_I�<��w?�-�=1�u>2�w>D��N�?;RL�g�>ǳn�D9z?�{8>�pJ>��7>�+����>�z�=o�t>#���|j?j8>D��=x�>yA�f�>Y٠=A/%>#ʠ��j?�Y�={>J3�>{��2�?���=_">*/��t�g?�K>��I>�&^>7�E�?�=�$:>����Y�?�3>)�_>*Jy>����d�>� �=��h>�5}?<>�ZO>*�{>�m	� �>��=W�=�U��D	z?8��=k<3>���>�>����>���<��*>��R<��?N�*>5�f>��f>��
�Z��>��=�q���_�?�uA��s;�5�?J?��e@?21ÿ\��J쭾�?�?b~]���1��(?<�@�GD?�+��*��<���ۢ?��g�<�D��9?
�2�-�6?�B�������m��+]�?�A�9=��'?~�2��'&?B�ǿP���������?,'Z���;���
?L�,�G�9?>�ѿ�R��������?�JW�� K��?�3!���&?�3ӿ�����ڬ��,�?�8\�z9��Y?�e�y\,?-ÿ����[�[�ٴ�?v\B���,��J	?f.�c�=?n�̿?������c��?j�]��r-�&?(�9�-oH?b$ƿ����ǖm�k�?x.N���Q�c?R�>���J?��ҿm������Q��?�'N��	9��5?�(�?+E?�ʿ����y�]�]�?l�N���N�U�?472��*J?����J���X�L��Ԗ?�PO�$04�a��>.4��zB?nͿׯ��]�l�+��?G���C���?.%�Q�.?�FϿn~����O�qÞ?��W� S?��<
?� )��p4?�Q��/%���ƞ�#q�?�Z�p�J�c� ?�2�WW'?R�ȿe��q���X,=cǂ>�|U�$�?��?򷿻C�>���>-h���e=��v>��8��?)�?�굿%U�>�0?>����F7=���=�]�2c?<;?_r���A�>��>����Q�� y>��[���?��?�C���T�>�ϟ>���P�=2�I>��8��a(?�?�?���1�>��>ug��L�h>[���?�^?o����e�>��>7�
���=4Pl>TeA�Z�?�W?������>��=>�x��� ��xL>��U��?�U%?c۶��9�>�u�>��þV=d^w>��P�^O?��?KѬ��Ĳ>�?>�F�(��غn>\0N����>j?ݻ����>�5�>ب����K>P�Z�`�?��?	Q���>Ok�>�����ڼ��=<Y�W�?��?����>[ީ>�G���<4>>��\��.?U?�ⰿM�>ݼ�>/����<B_O>6�C��W?�?G����>\�~>���S��$�>��Y��_?}"?����!�>wR>3�������}�>��5��7?Tu?�k��љ�>�>�ľW�x��0�?������?Гľ��轁 ��c�>�g޾��o�Yz�?hӀ?��Ҿ�m������>��ݾֳm��?W��Ń�?2
����9�����1�>g޾!f�qz�?'���x�?�6��y;`���W�>/eӾv�]�SV�?���K�?���74�x��-J�>�dʾ8�y�U�?�����t?�E��$ID��5�b��>Mt��o�w�	��?����}?�����7���)��>�\���'d����?�I���n?�۵�N.W�Q�ξ���>����;V�uݓ?ݐ��bgx?&Ʌ�ٷ޽�ܾ���>3hž0�v�h�?�Ӎ����?�&ž')�����5w�>Q}��_d�+d�?jv���˃?�x��z�<���پ_�>yھ/�e���?2���i? ���K��B�Ҿ�>�ƾ:�d�3��?�G���a�?Ć������@t�?���Ru��?���y�?����� ����r ?O����]�đ?�뛿�u?r���p�=�ɾg��>�����w��b�?�*��忉?Dˈ�5�l���G�>��w?�x�$��?�J$?�� ��?&��g�|�w6�?�	�?q*j��͞?��6?Xe*����?��:�i��i�?x�j?8}m��Û?�e:? �M��?r�=y���q�?Ngn?�"���
�?>�8?(W.�̻?�������g��?�?x ��-�?v�G?�-���?���]]����?�d?�j�����?([;?j%�s��?G�/<��C����?�(~?��l�6i�?��!?������?��|:��v��8�?rWt?�������?��>?0! ��J�?l��<@�����?z�f?H���R]�?>i'?�!��J�?�3=�*��c��?)�{?�$~�j��?��G?.�����?q�7�y����?�Є?��^��?��K?L'+��^�?�!ʽ[|��U�?�n? �js�?B�7?L?&�?��?Q颽:��cy�?Z�u?5�W���?QA?�p�S��?��U掾�?ͅ?LH�0�?ʁ8?�96�3��?*�{��h�s��?�c?��b8�?�2?R9��?V˽wy�cf�?q~�?�+�)�?�X=?z��eP�?p�<�˓��P�?/(?-�(�'?p�<��v�K3�<[$�?��K?�@�(�>�7�#a?޾��IH���u�=.}�?�gn?�@���>��T�>�*�=�(t�}�����?��b?�r@�3?������>Ⱥ�=�僿9�?����?#0^?��@mw?7�:�~?���=�fn���= ��?a�s?�\@� ?��:��?8V���m�8H)�9��?��t?a'	@���>�.-�}��>��=S<��("K=O�?Y�c?�@} ?5�'���?^>�Y��e4��
�?��W?�
@32�>]��?�\#=�t�X@�=���?Q�e?h	@��>��)�Q1?|1p��z����<�޸?��j?"�@���>�U$�P��>��o=T���t7��#!�?�UV?�4@�?��6���?��'=���[�=D�?�e?_@'�?�H1�ˑ ?,g�=� v�i��f�?�_P?�@)��>�B�E�?��|=�kp������?�e?M�@C�?�$�KZ?.;z��T��%��<;�?7�T?J'@�S?a����?�=c���w#�<���?'�U?%@55��C~?�&?)?6��>"�<�*d�@ �����=���)�?�B?�z ?
�><�8�w�G�웖�܍^>a��)�o?�'?�V�>P�>��3�ڸ`�������=������?�t9?@|	?��>XIH�`�������5>�� �q�]?�^?�=?:d�>��,��L����ʞG>%����f?<�#?���>:�>��9�6�g�@ ���o>>h����}?M(H?y�?�~�> O���H������ >�����;y?l�&?��?4��>��4�<,`�򜍿��/>��'��k?	 ?��?ؒ�>�>,��/X��4���)}>sD ���x?T�?9�?��>�<�\��i����q>�b,���k?�(?wq ?��n>*H0�
Q�9^���?}>^����n?�s9?K�?���>>/+���=������!�=�)���e?&RA?O�?e�>�/��l>��v��4��=mE6��_f?V�'?���>J�>O*���F�� ���^w>%�V̀?)�0?k�?�B�>�wO��K������ 	>Zٽ�D�?��%?�?g�>^&7�|_f�^��u��=>���}�G��'dm��-�>nl��!a�b[Ϳ;���8�޾���������R;�> ���� ��ȿ��⾁G��ǁ����@�ʪ?����o��>ſ���Rı�aڊ��Fؾ�L�h`?A���'A<�4sʿ	������������;��gN^��	?}���6:��Կe���$����줾e������!�?ڭ��'U"��7׿w�����Ӿi�����q�;��A?�:����/�V�ÿ!ҝ�(�־Ǽ�������x�?\��E����׿Pō�Pz��K%���z��g½l(?}���٠3���ǿU���$����������?p}��?}���I<)�F�Ͽ����^�>;u$����"��1?�Ԡ�T2�r�׿�����E�Aڔ�io����#�r��>$���!��pǿ�/����������Ӣ����:�?aZ��9�5�>0пs��t���o���[~߾��ٽ��>��ek=�~ Կ�L��֑۾�觾99־9E�|U?����s	���̿땿�Ϡ��_��'˦�c��Z?�U��ٽ=�V+ѿ�B��l">py?�T@bTo��M?۩ ?2Y��cr?��=?~�>��>�Z�?^�k��E?�l�>�8���s?�S6?�,>�?�r@Cf���?���>nU��Zp?��9?�c>�i?�1@f�y��F�>zI?�os��Xn?P?��2>�3�>`�@`Ld���>ZU�>h
�`�j?�(6? �+>$��>`@�9~��k?���>NC���?�=?�2A>W��>(]@-|�L�?4|?HB����? �.?��=`)�>�7@`f����>�?=�q�ͱ�?/�?>�>���>���?�Fj� y?�?�Ň��Z�?��!?R>���> �?��X����>��>��p���~?x�8?�u>`x?��@��y���?�M�>��X�v��?��,?�G[>��>c�@�o�Tz�>�>�>L���l?
9=?;d>��?S��?�	d����>|�>Ɯ��Ae?�L+?1�L>
?S��?��Z��?�:�>*|��Gx??��>i��>.^@�J\��c?�|?�,���o?o�?�>~�>�'�?J\��Y�>b�>.���o?%�?TQ	�^���XX�=S��Ӹ'?�5��r��������𾌓�KL��35�=�ݼ�@?i��2μ���	��׾�4�A���6�k;��/=��?�Ǿ�}��K��Ⱦ���(n����:��ƽ�� ?g�>/��D����վ���Ѧ����=O`;��,?�=��Dc���=�RMվ6��ގԾ��<䊄<�) ?=�׸���ʵ�z������ =�ڋ�Q�%?�b��`N���G�����륾��=�w?=�2?�z���A7�l��ƿ �~����a�=�=U�?_(���¿,�뾲LӾư�����]�Y=G����+?�ľ"�ĿG��Jھ���1Ҿ��=���sR?�՜�^!���Z�$��X	�~Vվ,�<�;�<�y?+#���a��[B�~�����ߍ��}�	=84='�?u���4�ÿ�u
��h��D��s����=�={n
?�.���¿<K�Mh��� ��f����S=w�E���?����J��V~
��
�r��}ξ=�=M��+q4?1@��V���f��,6�����?��?|]E��r���'���� ��s??���=cC�����>ي?��;�$���O������d(3?{�=�z��Q?���?��F��۲�iZ���W1��H?Y�>EG���g?'��?�P0������b���I�$4?�}J=�ž(t�>�?�P1��+z��������CE?a��=��ľ�)�>&��?�{>���!۫�����O?���=a-��#?Qi�?FG�NG��W���1� �+-?4��<wM���?� �?�B��������b��S?��-<?xҾ��? 6�?�I�v���E��3�cR?�:��׾�w�>�x�?x2��������,,-�V�K?І=�	�٭?:�|?�5�ܸ������/���aB?f~ >yP���.?we�?<�G�\���3\��fc�>?w��=I�Ͼk�>��?VzA��F���곿�G���/?�=�� �h?�߃?�I��3w��ԭ�Tqμ�qJ?�J<;ѿ�.?�H�?�6�pλ�kI���W��L?�?.=7V�f�	?i�?�H8��浾���r{0�f�T?U��=.xs�i !���2��A��>K�L�R!?��?2x���;}�7��H���	����>{b�i�?w??��v���u���-��$�v���*?_zW�D�?
?2���-��p!�d#�׭�Qb�>'P�3�?%` ?�Ӂ��Fp��(�p�����{[�>��k���?;�?�#���ą���&��"��9��]X�>Ku���(?�,?�{��"y��'�E�����>�{Q�w�?��?1'z�&�m�r�!,"�y[����>g�V��4?A�?:q��4�q�#E��g��Ǧ��2�>��g�U�$?o{?�Et�jq�����"w!�+�����>�$M�6?�?!N{��v������������>�am��-?a?B���&��S� ��P��:��Y��>#�]��?�H!?IU��	����y� ����s?��f��p?�C?B ���7��,�����V���>��c��j?��
?Ђ��ф�N��D������Y�>�Id���?� ?����fi���.�9�%�Sѣ����>��o��s!?;�>l���X��>���J6�=z��=��)ų?�"?)J��D�]^�>;G���>��J>�:6=`r�?��?=I�yU�k2�>W]������_>���2��?jB?��<���'����>���������=�\=�?��?rG��H%�y}�>mD���=��`>�7`�eʹ?�D?.8�Oo �-��>	���=��5>��c�Ƿ?�?O]O�� �C��>�H����<���=�/߼�I�?�	?�@������>߷������	f>�?�=|j�?�s?w�*�i��� ?CU�6�;�.>b��<�5�?��?G'I���a�>��(��A�=v(>�{�=l;�?c�?�b<��)�`d�>���ℯ=4~H>t��;�_�?��?E�K�����>7��7=f�>���U�?��
?�d<�e�	����>y�$������A>E�=�+�?�?++6�f�#�7�>�K���7=��4>�^�<�??�?��O�iI �xz�>��:��=��>�!�=ˢ�?ɒ?��:�u����>���$��<�8>����V��?W ?Q*�c9� F��]h>-[G�<z�>�R�N�v?r>R�T�/�<g�K�&�g>����.??���%�?�yu>��h��>!�`���1>@�|�3H�>/��#�?��>��M�O�=�M�<�V>ņ#��Q�>���SY?k�>,oZ���
>\Zm�D�Q>��U��a�>���Um?C�>�/�z�>�ZJ�bIW>�RK�=(�>�V�D��?u6`>:�&��?>��h�>�=>�� ���?���[wp?]��>
J���<H[b��	N>��z�^n	?c����g?w�>��=�e��=�pP�2+�>�Y�$�?�r��Zr?˚�>ʽ:�"=�`d��@,>�:q�DU?�9����?�=�>B	�����<`z\��2V>dom��o?&��g8�?�U>�n��[�w=B�k��y�>�W���.�>'Q���h?I��>��E��=��H�p��>w�.��1?C��o�?%�>�p�n��=��S�\Î>��\��f
?���{�v?��>�����=�OS��ߣ>������?�y�4�t?��>�y��}>Q�O�.�9>O�'��X�>��1mn?�kf>����M�=�@׾w40?sm���
��#I=��q�*v��腝>�&����K�?;����ĵ��P�<d�t���þ5%>�7%���վ��4?K£�Y�����삿F{��W-P>ɔ'��Ӿy&?)᭿�����R�<��}����>��>��e��i*0?'��3d������͞v���ھ��n>�D3�N� ��66?s��޺�S����z�L����]B>�k6��5޾��1?���-���%a��ttt��~����>�08��{ ���$?i����[�ʈ��a�Ђ��Jo�>y��	~
���?�ޟ�󱍾q�Խ�^�~d����>ͭ0��\ξ]%+?qo���R���D���b�~�ʾ�9>-���;�/%4?}i�����d��< ˂�������2>�v"������%?娬�����Z�?��w\�,�¾ڐ>�J �.��U�"?��Yǭ���:�w�02оh)�>�8���C�?v���Z�؛��o������m�.>K�$�@��?�-���P��=��+}s���þ�>Q>�%��
���p?����e՟�Hb��gu��IȾ�*�>�L6��9ҿ	1���(?/r��c&=��[�?���c�ھA���W�ӿ<���Xy,?������/�,6�?w��w̾�T=�W׿7�,�B?����9J�\ś?�a��}��+���%տ��n�D�?������F����?۱���־�?e��Ŀ�%��E?q���G�1���?��	vھ��q��+ӿ�DP�l-?=���.�$�Y�?������U���Ͽ�6n�@R(?k���8*����?Ԯܽ#�1+Z<u1׿T'�2�;?�͑���:� ��?����Ǿ�_j�koɿ7�� �"?I⓿V�9�F��?�+-=��	�9
ν�9οC�7��1?����qJ����?Y����U�_}���-˿
Kq��Z-?k���VBD�tȎ?^ӽ0����%=�hҿдZ���$?K[���0����?V���S��Rн	�ӿ��&�b�:?����i4M���? [:��,���Z_=Ӥɿ��*�0E?񈜿��+���?.K���6���H�<�ٿ#�v��e?u+��U).�$3�?�ν�
���ƽY�ǿ/�K�P�B?2���r)��?��m��T־f��CL����u���?V��<�1^?~�u>��a��w�K��{+��l��p�?Kڂ=�7?J�y>i�p��O	�?���KA�Ÿ�f?1=�A?�5�=��j�� ��D��#c�Șƿ��?'�����E?6�j>8�G�UJ��Oi!��?�Fÿ
��>����[�@?�+:>��_��1"�!�9�����ſV>�>l�J���U?GW�>��]���ٽ�	�����R��� H?�B�<��H?F��=T:b�e������/�bT�����>�@K�%CT?�=>�NU�����]�q�������?3Ĵ��*E?�~>äk��ȿ��,���,��'ƿ�?d����>?��Q>S��;�gH ��g���ߒ?)����C?Fx>D�L�S���Ş�͹��0=Ŀ� ?��k���[?�$> _P������o�=��,�>0z=�T?�]o>ռ\���x�1�M�>�(����?Ӄ;��O?b'9>�c���!�����G�hǿ7�?0��<��E?��>��Z�"O�������z���@��>�<u4L?6wz>� O��q�%!��𸐿yQ�=����م?[]!����>9���U�n��������=�	��?�K�$,>덄���c<�-�ㄿ���=9.��=�?�-/�n�V>�󁿴H�;d_G���}�/=	>�x����?��?��>�az��s��ĵƽAe{�	�<=T��?��ٽ�8;>.G���*���F<����?�%>?�!�N��?��ݽ"�<>Ք�ﱙ�I�(�`��u�>z�����?�{ͽ��>7�z��}M�-3�^߁�->� ��,�?XC���d>���@��8���{��� >�~���?�+��9>Mv�lnd�#�k��n��Y >�y�ˇ?_7E�:�->�4��d�:��1��=��i.=�T�Jb�?����>>��s��򫽋�'�������9>�����?;^�S�>�B���9)��|���쎿o��<�.2��%�?�*�b%>8[��K��,	��t��7�=s���M�?*��P�>ә��e�%���н ���+�>�[�>Ƈ?�
ҽ8t!>�U��זս�8��凉�i�_=�%���?�����\>����z��Z�>�+;��r?'�>��\?�S@Ns�=�D��s6�;{�J>Y�-�#�k?pN�>;^?�i@=0h<��j���<!@>e�9�y�`?�=�>�~_?Y�@�� =qԨ���3���>5���xj?I�>�Q?�y	@���=��T����u�|>�&.��BO?ʂ�>`H?�x@b�=}邾�P�<õb>QZ!�1Uk?q�>ixV?��@n(�=}�>�-�<I�q>=/��so?�y�>a�T?Ԙ	@l��=-�X�kf�녓>?�;��j?���>7�a?@=@a�,=�ؖ��V?����>-���c?Y�>�Sh?�z@��=Y���}�=;�>&>os%��U?HE�>��P?�*@k�=�>���&=GS>�';��oq?�>�>�l?��@���=��c�J�*��W#>���Od[?���>)�Q?Ş@ ��=/�����==o}>�c'�W�l?�`�>�wV?J�@��
<Ņq�c�J=�ɗ>�)�[4P?��>�e[?�_@���;51U��)�=���>;S%�&W?�ԏ>��c?Y@Mx��B)���#�F4>s{=�k?M�>�S?��@�l�=�u��$�=3��<sJ�:�|����?����O�@��Q?q{T��]*?��c�ݬ�	��<���?�󉾹�
@8-_?0���!?9G~<?K���E�<H�y?�p�&�@R~a?C?ҽ2"?o��:!����wb<)�s?k�R���@��M?L�=�N?#5нIY⽿(����p?��l���@N�Y?ɭ�;��3?<&��˿���[=L>�?~��l@��C?B��
�/?A%߼j�ѽ�|���?%�j���@�\K?	���6?<ۛ��>��%��<��?@��5�@�F?�[Ӽ��3?��<�H��D���S�?�B��u@�Y?���$>"?z�<E���?ۉ�/�?�3�C�@`�b?\�&=��(?;�eU���Ċ���?�*P���
@8-]?YX��v?�V=�����+���s?�!�.8@��\?�==�?x2><Vxb�U�=B?r?�D�RK	@�@>?��+<�^?�xO�O.��چ�Ǘ�?f�ag@&$H?����;!?�5�f����½�΄?�V^��x@D_C?I��;� ?Ћ����<2^��0z�?����D@\'Y?Ϧ���V-?�,?��>���f��?$�>m��`�X�>8�L�D�.?��>�~��P��?Z�>v����T� ��>���ƀ,?��>�v��п?>d�>�\��pW�|�>*(��0:?y��>������?�bj>�B��sg��6�>1��<�gI?i�>"!���?dϬ>����Ii�@Ř>e.��_>?�P�>I����?��>����?�Z����>�m<BB?��>�4��(�?d�>��	M���>�H���86?�>Gt�f0�?�Vk>���[���>kI�<(??��>��ܪ�?�&i>y���zg��Ÿ>Y��<,�+?/��>����*>�?��>2���j��M�>ȖD���B?[ӷ>d3�>�?8��>A��s�d���>�c&=��7?�n�>�I�,��?f��>Y7����V�١�>~�m��Y??
��>Dv�V;? D�>�ړ��
l����>�ѽ�>?+�>g�N+�?�	�>��˾�b���>��7<��I?߈|>�� n�?¥>�ʚ��)O���>f!���W)?���>�G�?�px>�J���Ag�O>j؍�L�@@�K=}%�/���sqj�A)>��>��v��
���@�����?�;ǳ�K�_���->=Ф>b������� �
@>n=xO����yHU�� �>�ʽ>�1��^��҈@f�0=gI����]�=�(>u
�>d��cg����@��,=��#������U���H>�ٹ>�7�����&@�^G<�"�Im�W�I�cu>!��>	����匿:x@W�<��*�'�ƾy�m��_%>�ܸ>�Ný�Y��dt@����%����k��M>�3�>JC(����
@�β�o�"�� ʾ�4g�F�k>6H�>8[f�c����p@7*��J�"�Y�ƾ�i��D>��>7�������m	@�ƽ#2�s1��7�l��I>�Ʒ>0�i�T�����@\���{��訾�"h��iL>���>[�ͽYe����@@ύ�x������6c�Į[>�f�>�#�*B��"�
@�G�� �����+vP��%�=�>���x��ȸ@�2<��u�������[��>t)�>���)��dV@'j�<6��h�־��T����=�>�9�63��x�*>h��?m-�a��z's>���<t0���5�>{�ӾBM;>(��?��働��x�>�����Z��~��>��߾1d>ꐇ?;{��`���M>�|z�P�׾�f�>�h �Á*>�?�k���g��Ҏ>%��.r���u�>�N���Gt>�=�?����\�+D�> ����K��R��>�3̾�>>]�?�y�Km����|>d�E��N�>�bȾ��W>�f|?:q��j����i>��\��Ꜿd��>���,|>��?���P�_2�>o]����پ@��>aȾ�Le>�d}?V�g�����d>	d�<|Aξ,�>_����>>4߅?0��񈥾r�`>,�������L�>�׾&>V��?����DY�S8�>��� �ξ��>O�S1>8��?M��-����>�vĽƭ���>>޾�>�0�?����m��w��>|�Ľ`�ξH�>��۾6�=>!�?aY��:���ǧ>���
砾��>�nؾpʌ> ��?
��}NX�錂>
���Pپ>,�>��ɾHWe>C҄?e���%���aS> �½챧���>I���8�>�̯�	�������4?6�-?6��?�?����2��>'	��B2��7_ξ�?�.E?�@�?v?����^�>�ȱ�����nf��!?p�,?�Y�?�2?Q���3�>E��D夿�ľ��&?v#=?�&�?�]	?���2��>�[���R���ʾ�&?��!?Z_�?ng
?���lO�>9̫��$��}+���7(?�<?�B�?���>���� �>E߬�l�������"!?��#?
��?��!?U䷿4��>/��F8�����m+?l�'?�ڷ?�?�«����>u���������-�$?�e8?XS�?�-?���ԝ>-婿:,��S����?b/?T�?з?�׷����>����j��c)žM�?R�?Jl�?���>1[��(D�>Ϯ���<��� �ņ4?:�9?�s�?^	?ù�"��>Ot���Ѳ���)e?� "?5�?�?#����>��������O��˧!?pb ?4��?&�?{h���Ʋ>�ϭ���e�̾��5?(�)?�T�?�B?�E���o�>%#��xr������5�/?��2?�9�?��>aA���9����>uڬ?K���9q?��A����91��2E?�r���=Y��?SX����v?�N"��x��R�!=�?2f�ܸ >c��?��̾Bu?'������o�<u� ?�pw�-V�=]!�?�ɻ���|?�94��@��,(g=�?Xr�|�<�+�?+Պ��;�?4$�*⬿r��=��>��g��{p=?��?h����t?2�2�Y��?��=�7?F�}��*]=�K�?8����w?>q6�L���A���?#Bt���=�p�?h��&,s?��%��F��"R=��?6ys��=���?�u���d?�]�D|���F�=w ?�U��[�<��?Dg���n?59�ϫ��E�=�?�瀿G��=�b�?�k־C3d?��!��*����=�g
?zL��`�=���?�/��)�?��4�v��0�,=B�?�De��r�<���?�9��xl?Ԧ"������T�=�L?����y�;�a�?a����k?^�#��ʳ�E�=\?x������=׺?vV����y?�,��L�����;�?�p�`>�ʹ?����kwt?�<4��ֲ�05U��	?PKIVRN �   �  PK                      archive/data/1FB  �
�>���>G�=x^��B�>*j>�K~�y��[(����R?G�4>q�>�O���������?�� ?�x=#?�� �Q��a@ֽU�G������>[v��Ͼ��
�ͽ0S@z.���>�~�~W=�e���W?JgS?�?���.v���Q��ِ�:0�h�>�Bw�ӝ�?�n��%��=�ї?�:?�↾0Z�>��%?D�>�G�u�H?�[<p!?\�������b?;���b����2����PK.��      PK                     C archive/data/10FB? ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ,�@���@Gt�@�S�@PK��)o      PK                     4 archive/data/2FB0 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�e	@<�=�$�@�]�>	f@+�@���?C��@E-@�[�?8�y?4��@(\@�@��i@��?�?@̆�?�B6@(+ @�s�?�?^F@6�?1��?��6@�fM@Z��>�?�51@74@�Ef@�R|@�=�?
�,@�K�?�x?��#@�r;@�+=@�[K@Y<@';?�{#@��?�E?���?a��?^J@Hf�>q�?l�1?%��?��J@�Ǒ?�k.?�Ύ?�'@ע�? }�?� @���>9%f@H�7@PK�PX      PK                      archive/data/3FB  ��@�������+�?M?ç��rD�ݣ@T� @ͯ�?x'�?�G����#?;й;3?;>3?Y����?N����^=<l>_Ȭ��Ζ?����H���ܮ�k��[9����B?HY�U~��?>�Y?9�>U��?o��>��?��,=HL?�?sM�>Mj��9��?e��?����ڗ�>6	��~Y��}��nQ���=�?S�F?D�K����
@�H�?�h�?"'�?���E�-?%Y�?�]�?̀R>PKv�@�      PK                      archive/data/4FB  ��?g�&@Xs��]UA�"@X&4A�A�9�½����'ݾ��T�I� ԡ@�A֓A�������@HuA�.`@�e����.�#I,A���Wk�@��/�b���R|AP2A5Y���S���@@g"�/�M�)������@�!��v"A��@oL%>�>��0ʤ��d�T�$A�D	A�����J��%:A' ����B8�N@�������@����Do��BJ���Atc"A��@���*l��	�NG1�PK
��      PK                      archive/data/5FB  2�A�d;A�JKB\�yB#�B�f�B;�B��B�%B�B4��B�^Bx�(B~1EBQ	B� B���B-�tBѷRB�R�AU��A� BkFBڛB*�YB���A�C�A��A;cB3��A�&UBPo+B�RQB�$2Bx�B�CWBR�YB��]B0�B�BMr7B�K�B���AE�qB��B��Bc;TB�3tB)�JB�|�A$;B�1cA���A�m�A�dB�o�A�>A
Q9Bj�+B���AuNBB�A�|hBѥ-BPK����      PK                      archive/data/6FB  �x)     PKY��      PK                     < archive/data/7FB8 ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ�r�=d`	>d ���j����>1���3�;=��;��>�$��]W���3/�>Pe��R���,�>����>�����>�^,��h>`��=�c?.�>���K�LV�>�#>a��>,!
>8�>�;�˸�>�W'��v�j�>
}�=��4?�����Nc��\=؝�>B�E�,�����+�ž�7:>K>Y�`�Ī�>81�>�t��K =�h%>�6 >�)"��]�_�Լ��.>NKڽ̾M������DI>�､"*�>��G�� =������>�1G�����wƽv�>��8���վ�
��R��>��;=�
>�80��`?EL>\x����o�>h���l@M��;󺭚�>�X��V痾gկ���L�	�@>Y�=�c;<[&������q>�r ?X^��0��r>�l�>]6]���.���D���P���x��gt >A�ӾA.v����>+e$����G��!��>*Yü�O�ٺ��7%?c��>��
=�����m2>�/>���<�ꕽ���>gٹ�(Vl�H0]�jө>=�н�"۾T�Ӿ !�>���>.�C=�'h��	�<#D>Y|�>; ��t�������> 
��	7���G>�v=d{��nt��e�O�5��D�a!�=�î=佤��hO�>��>uN����!�3:+��u?�:�rӾ�����[T?Q��>{���FO�5,V��Wj�*@�e���j����}�>P�{>m�\>������p�J��>��=3����[)Ǿ	$��8��>__>۷�����>�f�>;���2`+��K�>��->~A���׾.��=�K>�����H7��[�<Ғ�=#�`>��.=
W/?GI�>*n���Ƚ����=F�`�B��\��p>ke�=�+��B������#�����=�>>]^?'>BG���z�?S>f�I>\ǀ����+��=O�>��>h�>�pU>�'>�IF��%�����C<<Nv�>��*>�Ǿ�Z�>����X��>��}�8��(���X��i����0�| �j��i�>����~��>9-=�By>=����ܷ<j �>N��>��'�����6X=�m�>��>�����,�ʾ��;� �#��=�b����>���)�*�F�*->���=M�޽�帽ma>�)�=
�)=g�o>���>fU>Y;>�-?����|>��>��>6;��\v�;33�=�kV�(���;���q���w$���>уR�Uj��1���n��>�1���Ǿ�����u�>�$�=��%�5=>�g�>Cо.�T����=sl־to�}^6=��>Z��S(I����>0��=+�+���wDQ>��<C���<D��v�_��;��e�z�mJ�>�+L>�!*��0l�j>�_�>�����c�K������%�|��=E3<e}�����>�$e>�T��9w��Z�>oҥ>��(�����,>���>�+�>ͷ�>�Z�>�{�>���JQ��Hi��%*Ľ���>��=��>ϑD>��H>p�>��<b�g;@ �>AN�>�u�=�M�c�J��>If>W�����m>	#�=z�=�þ_�\<Ԡ�>��>��R���־.�>F��>]LǽAA���� >��ҾSY��5%>���6?�H�>xo��'���S��>�w�>�	�>��>���>h��>p~�=M�j���������l��>c5�=wT!>I�n��`��i.(>���>�hp����y��Y���ƾjP=���>M�=�����O�>Kw�=�'��v����#L>]�>��6>󫮾�j�
�
>�>Aa>�g>8<D����=7$u>t:��C&�L�*>�=�>��x��a���O���0�>$T�;�� �n�=T��=�b>\!K>>��(�>¤�>�?ҕ߾X��>��>���>"�ݾ)�<�!��p�F�־V!d�������6>�@��H/�
z�=��>�ӗ����Y��>�L>Wi�7Sɽmgi>,��>��=�� >eg��0B�>sx�>�#��ud�(�F��:�>&���^�-��]��M��>�h=����<,��>e�/?�Ja=�%�!3
��5R��e">#0�>�k侘�>��=J&���c�eo�>p�>:�$>Ғ%�}7����L�=�tu�͛E�&>&vc=i����v����>�H�
Ë��6��C�>2t�>x�>��>��>nCv��:�>�?�>�v�O�>�����ӫ�πd=��T>�n������w��\s�^I����>��=���>��I�[��>��1�/�N=����w�<>�k?�Ⱦسľ8>=?�7�>�
�=�=�ɽv(G� P4�h�\<�:�>��>���Z��=Fw����>�p��䜾�5��8�;����]>��>J��=��1?[�=�}/��/�={?�X">�\�����T��>���=�̎="M^=��:>��>�$a>�
���K>�٘>@�f�`��1Qu>v� >�Dn��cϾ�=%0>�>ͽ�'	��p���>�5u=�d'>���<��v�\�<�d�=(�Ὥ3��F=_��B����I������A��E�>�>�FT>uҾ8M=��� >���=5v�	�>�
�Z��=�_�E<�D��Xg��f�a`�����:=9j�>��ž�>�E�=Θ]>�ž���=�	?�x?O;���n�F��=m�?9pN>�/U�_�X�>m���
�*��>.��>�f���u��(���>�&���m��ξ�\�/�۾� >#��<K��T�7?
�=!���l>�O��>��X>T���sѾ7�>jO\=�C��F�=M�S>@>�S�^�ٽ�?`i?~�����<��>\�T��̫�����Y7>,��A�>���>�!�F��>�~�5�[?_�?�H=�[o�=�l�>>s@'=b�;�FF<<!���m�d�$�#gv>j��>��>�N=ݿ���j>��N=��><��YUC�E1>��>��ܾw�ǽ�k����þ�o����=�I��cIҽ�%�>._�齶={�C�W<?Z��u����H>�`N?�����@����\�>&o0��y�>�N���Z����>��=��?OU��{&�V~=c�>���� B¼�_�1���H>��Y����f���>V��=�|��ů>b�y=�4Q�9���z�x>�b�>���=ܲ��#�1<L�/>�Q>L�\�A����=���eW�ʱ�=N|�>nر�V^X�켟>��>Z+��0U�荄� :�<�B�~��>��>6��������>�¾�*���� =��>y�t����h���>�í�M�������.3�6����=�m�D�߾�@�>���&\����d� >�H>���r�~�aG7>6Y�>�d&>kdu�q��2��>9��K���߰>��>�u˾c���8��>4�>+7>�����{b>�=��Y;B�ܾ#��|D	>�i*>8Y˾���>�K�>BR>Tо]`�>SZ?Os�>R� ��VH���Q=n~+=h��>4�3>�}������ �>��оmj����=Z!�>w�9���p-����>�{4=�&F�����>ޞx>Ζ�����?>XѾ�H=���>
	�$�
���-�o��>b&�������M ���ɽ����2��>m��³ռYL��C�>FL�=o�\�<�E�U(�>U�'���A.��%�>$j>�!@>�#��7�����>ˆ��OPԾ̷��'�>�1��i�&�U��¦>p7>X����s��	p<ASK?���=�|?F�,?��� k�<3��<r��=�*�;�4�m\�=���>��P>Er>)����~>@~�=b^>�ʚ�&�>�D��&��g�_�ԡ�>}�D>𝾼��v�B?�LK>�0Ƚ*����>��=ڝ�������ެ>����E�л����p�>�Sʽ���
��2/?�>�(�1^C���=�[��G���GȾX���NP]<��1>J3�x�>�>{<H�ռ���?1�4?H�A>ɴ��˾"�ڽ�C�=h��>P��=�Sܽ ��an�>�آ���=r��>ҷM�����KT3?ʌ�=��=�_����=5b��,��=Hݽ�ѽ%Pc���ɶ��?�c�<ad��2���An���=2��=-s�="�=�+�<�mF=^U=I��<{��<_�<Jړ=���<�5><d�=��>k�=ţ=O�=P�>u^w<h	=�(a<��=��; w��`�μ�>�=*��P�P/��C|���k��5>S��=�2]<�>cCW=��üB,R�F��q<E����=���=�=�g���
ȽG�3<��<��<��9�|=�=(=<O��Q=���='���}o��]8105>�]��X!o��e��Q�=3{1>w��=�?�=�=$>qɽtw���6=Dʚ=\X���_�C�<W@�="@=�
�#=���=N~ϼ ��=5���<&��<z,�<�y�=��]=���sl=]��=�@�����)�
��ҽ-B̽I�=js�J"�����-���D�<F�ʽҰ&��'�=(~�<'�<��(��=��=�9l=��ٽ�"[='��<F5��!=��=#2=����=��W2�=ȟ<��ʼ����u�z>7�=q�<.��W�7������5�'��O<S��=�e�/併������ ��a�с��Ə-==&��M��G�=��ؼ<��<����5N�=M�����.������)����4�>���;}��Gļ��½CN����m!}:���>���0��=e��<o���`�j<i ��ˁ�;o�P��䓽���=��M>�C=�4�;�S>��{=�Ƞ�s�����X�*tk=�T��;9��#&�'�=�s���$X�S �<�[V<t�g���=E�$>,�>Q�G�\+_��Ϣ=p~9������=�S�;��Y�#����s�%H���=�ދ��;>0;�=�`W=VT�3��&��j��<���I����v�;�D&>u��=�>=H��=�7�=��<̓.=JZ]<�+h=���&��p�;�r�<(Ƙ<?=H�^��|��`d���9��>������¥/=��4���y<�)��{�;(��=���=U�[���(<�ƻ���=C���ٛ�3�=�]�<X/ɼ=᪽�fW�*D�9�C=��uɞ�	?(=t��<|�=�X:[%ۻP��4F`�ay�=��=��=!\=՘=G�3�;�[�=�N��~_����)<�Ύ=I�<g3�ȗ�����<i�Ǽ����m"�=[wD;�����Q>�W������'㙼r�=#�׽�T����׺�>�#�=���=�J>o/">��}<���^����;ҽD���P<���z`������NH=�a�<a�P�_(&��Ҥ� �:��?�46��q����V��b��[ =�p�=�r������i�<�#<����-�0����3�<M��r��=&��˂+��>H�=�g��24��ʎV<0~g��)�
�<�z>8s&>v�s=�(�=�q/�?ⷼ1V*�du��
����= �H=2Ӽaj⼄��;�=�=��=��b<��=�"�=8h0<D�����=b<��='��|5<�K�=C�>�47����.��i!>��*�<��<�==�=uZ�ʢ����ü^�0=9���4 o=���=�q��B�	j�;�d>=�)�<��>�`�=���=
�d<��=y�/>� P=�P>GT{=cP�9*`b�]�$>e%>��㸚9�<%[A=�	_=�f�ɷ�<�ȗ������=UX<E͐=!��D�=X2==��=2���|��=�M�=��q=)aýf	�;髈=3+=/S>��������=��=Ѓ`�H�-����r=����؍<q�ļc��=�qC<!d�������ǽ���=6 ���e���T;�BF=�D�=�-A�=աV<��=C��lL�/a����1<�� ������e��0�^�!�g�R<x
�<�ּ��<ۣR=+,�����T
�"6=ґ&=t񀽴�N=&K�Ӡ:� �U>������qeؽ�5�=�����̽s����=���6�j��Z�<� >��=gK���Ƚi2��\e=:(�=������z>k�q=2"<z��@z=��B={-����N�ӕ��xP�)�ӽ�$����=���<�2)�mC��s�K=V�d=��V;����n�Wm<�����9Ͻ!=$r\<[)ǽӻ=Y���;A����~�:o�N=\Ub�FY��#]��U��j	}=I��Wh�<��5�4'%��jٽ��,>�r�;�R%������B=:�y��D��
�L�=m�<J8������%��zb<Ҧ�%��B��.�=>aJ��ź�Or�<j2E=�?����e��� ���� 	��z�>#�)=m�ټMa>�(�=�a�F�=A��<C�5�\3��N��R�>���=7�;T͝<���="�=7�D=D_�<�8�=��=��ѻ�F��4=01=>f���ǼP���f�=�����ܽ���Qa/=�޵=�i�=�m�=$�=�}�f|;�<�=`-
=�ҽ�.�<C`
=e<��+���G��3c=}ػ�p��=��� �-��)�=�7�="�=]N�w��=RĬ<�~3=�\����]9삼O��;�3;�D�
�&�=%��o=77L���ԼQ��=7��=0��=I�<)�n=]��=#��P�߼kĸ=d�s=�}d�*FC=�ҽ�� �� =T+��ժ��z�&=���%:�=V�=Y�9=��˽�B��@L��%�����=M��T�>i,�=Q9%<��ʽ,��<�w�=;������a�H���<Ui]=�O�:�=�w>&�u]=ݭ��ؒx=Po==?&H�l��t�<9-�=I�͹��xT=�5�=T�=�� >��=$z�<�J�=ҩ�=���=Ԃ��
�=H�>+T����V;�b�]>=#�<���;,@��{����-�QG%=~�=ei��5_3�p��;��=N�����}�=��j�.4��A�2�˪�<��<ES���x��=��=��7=�	>�1<�W�o��=��>�WȽ!}�<�]X<��>I�@�G¼?�%�b�<"g;�NI�=�>�!�=C���G��=yy��_sļ��g:[�C=\�=���q�ּ�i�<��ɽ�<�l` ��!�< �I;΄�;���O�<���=��=0B�;ڎ`=�<�=��=�×�n�=[c�=�i=�y ��۾=���r*w�E���g	�=��0<c��;v��;���=!ӝ<�Tͼ�����l����<S+�=�瞼�����D<��=��J�����j潷k=0�8ҽ�bн���=:� ��B��SCO��֍��P�&���q��S�S=4��t=~w��7p<疺)齧�м�6���<۷6����͚.<Y�(=�,�b�����=vnl��񉼚FD=ӵ�=�X�;�c뽬���9O=�j�=*d�;璢�j�=����
5C=����y&J�?1P=� >�R5�5=�̓=��==I!��Q��'�^<��;"�=ubq�k/!�e9ҽ���=io�8���$P���t�< �L�m���@�P=��p�����_���=�|�;��㽇o��pЕ=.hY��9�Y�ѽ�,�;�4%�|>���5�����=q�t���-�޼
U=G���i���A>
����R:?����>�H���N�ߞ�K�y=㯽��⼾��<�R>�>�����WE���V�SA�=B���Fq�#q�=� ^�=���)y��)M�=1�=F	���ṕ=V�����>���=��=�E�;	�=A�=M�=/��<W�}�=J�<�6 >T-�=v��Q�=�-�=�X=���<�~��I�=\�&��j=������=ZY�<У�w1W�h�=�[�<�ꪽ�����H�o�0�T=��sؽ��<�K��������Q��)��r���L	�L��=^���"x��k����=�oĽ^��ｰ_�<���<�f��;�K 6�4��<��=S �Zi�=��Y=�h�<I[�<t�c��̠=f-���4�=�ܰ�o��<9.;'��=���Ŝ���<�Ӽ=��t����;���=k��>�O%���z�]��>��C��O���Kٽ�X��u=#���~l���V���=2}�z�a���>�:ž�?0�?P�>?E��>�$"?c3=��%?}�=?!D�>?T�=�P$?�K^?@X=?W� �;��>�:�>C��?T�_?��#>���{B�,�!?ɴ>a�>ճ6>z�-?2.��>����!�>�������a?ˍD��(|�h�?�r�#�%��P�iˀ>*����%��s��0��FD-�{��>�E'�1c?�?k(U?}��<?��ؾ�Ng�W�j>��>o��p���(w�]Q>D�w��({>X�`>z΃�r�?��?�G�=Ȗ?�w�>��?>|N'=3�/?((�=b|۾�}P���?�K.���h?�w\�}K�?�#�o�?+?Oﾪržj0E�1n�>w�_��_����x>��[?�6�É����U��5�>m��pV/>�g����K�=H��5>Y�.{�������jt?,56=�l�i����5[?��>��"c?V?�7��Tž��Ѿբ�>�ÿ�|�r/>���>E�+��Ϝ��b=Q�>D �����=�@'>����#��p���i��<�=<��\����Ѿm$�F{�>�Ă>.���!+������>�i�(b��n��@�� �=��>���MB���AɼD�Z?J[1�Y�8���\�B?��2�@#�0V?�ǈ�B��?�.�>�v*�"�ƾϬ6?펄>�j�=��=��>�D`�x�=׮ѾT����<Tdd�P�>2�ý�-��T�r?=k>Y������W0�>���=��n�ݒ�df��O���>�[��*<?��(?�ţ>JUu>v�[?bլ��Ǧ��^�H�`>������V����Xr>��F���F<��ｐ�#?��=��>᾿8?��># ���t]��)>m$>-�9�Y%8�i�m<�g�='�,�Ku�!B?�?��g�䔻>gb�>&��������mt>�'����>XY���f��ğ�oZ־�n�>Á ���R���E���v?�1?av軀cо�h5?V f=�	>��O�U �>��R?�*G=u���#
>��>�w���܊:��<O��@���o�`���h��ν�_�>�X�kR��Un>̐>b�=\
�;]�?����,�0��h��z�>��2��S�>Q!�>VO �H���s�=}K>x�?е�WP?��$���>��4��3=`ܡ>�c���A5?p�x�K/>7�W=D��>�����>P�O�@�)?!L3�OЦ?Z�@�G;'?�_�����;3�>�b�-������>t<��4�"�G>8�M>rc�?&���>g(۾-��=���O设��>HF�/7j�$���ɪ�>���> �P��q�Jju>���>Y1�+x�����ߑu>n�u�~�y��K.��^�u g>ϱ>�z���ā���>��>�o
>�C.����=y̆>�բ>���<��?t��[��
)�	�?�;?@��>x��0$ؽsC?y�+?��U>�П����>;�g>:W�
��<i�;�|j?*�>�"�<y<�.��>���>&>�0,��G�>�?k@�>�<|��>l��>�����"��5B��G��Тþ����EP(?s���,>'��>u�K?��w?��Q?��]?�\������E��8�>�  ?��Z?g�	?��$>H'H>�a�(�>(��,�~�$�rR/>d`�=����A?��
����|�>#�V���j��e�o��?��~?��9>�兽���>��J?��W=��2����>["r?����x'��1ݾI�4>�Y�>�W�>m�^�(���d=��\>�3��TX��j��� �=�U�]2վZ�?'�)�nlI=�eO>�"����>=�׼�ͤ>�]�X�N?��վ�y?P��a�=bIQ�]>���|S�� 5�?�1Zy����Zrg>��=�t3��{=�
?z�?:s\�$���!���?�Q�@�뽇2��A���'�>���=�>����޽�V2�2����I ����><Ǟ�xK>_����1A?�4���uS�yYh�t�f��
ŷ�}EE>ܧ�?�>YiC>�C?�h��F�=.@�R�?����.���ǌ�6=�z���^ȾhZ����<:�����kf6?�zR?3z$�KM��9��I�?���f�>��>4,O�#���L5�=s����m>+F�=�>x�[>�3�Z Խx�e���j�� �U��Z�>�")�Z8�?l�<S��>в׾�̺�:˱z>��0�4���6��?�1�;�� �!�?8�>�y<8��eg�Q۾������Z�����>Yp쾷�'�dJ��.����iɾ�[����m(�B��=�"�>0�?��=>oU|������B:? %���j����R�l-�>~�%>���)7%����>��*?��c�XU<=�g?䢙=YIP�v���R->�0�=��v1����m��]�<W*f>�tk�}BT?˪�?x�I?��&?��?㣊�L�>�w���W>Hy����n��ܢ>�?�=nQP�P>��\�nOw��'>o�>� ?qg��o�>V�T;uO7������>?�"r�3�d?�h|��Ƚ�8[�,>�]'��'�W��?��ȼ9�:��+���"?��@?�8x>Q��F��>��?�M
>��X��?�*#?o���#Th?}_8=�Z|>/�>6G���j8��~>6>�0�>C��de#�D_���`~�7�>��A��>O�<2c3;�?��D?���>Y����ʾ��I?��F<92��J���E�=� ὜Ҿ>��$��=D>?ͧ3���0���?�?/?TG>�mQ>��>���>�߾�l��o?l�O=�Е??V��ޔ?`���&�@?�6������r&?�Xډ='q8>���?�ʽ/��=�e?��>s���q�>ֽ�>ꭐ>��>��ܾ��>�'���>>9���Z����z�e�� +޾�Ὰ ��K�>B����><)^?v��=��>����+F�<���>�)�>N�=�z��VO�>��>7���R?7�ž�i�tU?,�]?sh?�>� Q�B�B�X?�����M�>t�d>~�{>u9����l�K��]a>�˼=G̽G�>"%?��X���WM��]u?��Z?m�>��:���>��,?�U��N�����>=�x?Nt��G�;���
F�>g�V��pѾ?jъ>�鬾���a�=�f�?#IC>���>z�ڽ�`3?<��k�>5[�}�>!�?3��>��e��@��A��>\׭���9�l���  >��s`��e�?�Ce���M����=��^w�'�m�*S�U�j�&��y����3?y)�f��=�?d��?3B��*Ϗ� �4�転����W=��?<К>(�0���=1�~��қ?��b�/�>�Eӽd2O?����WnU?I"a=<�"{b�f��?*�'>�̞��8���>ق�?!|=t�o�>�ѽj�2-=��ؾ�r=0p�>
#`>����Ҵg���>�U䈻*ދ��i-��`ƻF.[=m�����m�?�H�>��$R�>�g?I?�>�o>�ƒپO5��i�P����^0��#�ý�ؓ>�	C�^^���n?|N����<����$?%�S+>CI:�e�>z2>`�3�
LѾ�&?j�&���?�[�s7?g����J��%ľ�@�=�J=?~X�5����>E66>�m��]���� >=a>�U�K���,�>U�3�" ?�7�>�iR?l�@?Ŝ��K��>�t]���h�����g4>�T>�?�>���������>��>T���ƺ<#��>���>��*��
�&ʾz�>5���J�j>�w��8b<T���|_�~�
>֚�>EBP���Q�DҔ>qO����>��6'̾k�;>�߽�ၿ�x��l,��SV�0��Y�Z>�h*�Q���.}����@�?8�����T��D��cd?tQ|>���>��@=�+y?�8�0�?bQt��<<���?I�>{�ys�I�>�9�>j���f�����>����}>h�ϿA��>�e�ь�>)�?:[<�=�<�u">�X>�l>�䂾����^?)r=&~�\硽��:�i�W�t/�?�Z��(��x��=��a>hPj>
b?��>� ?8>)	�>��5>QX�>z��>���=o��=g�f�.,ʾ����eQ>x������=q��>�<A�,�02>ٳ{?��>|��>��O�u�۾Q�n��4�s�>ʄJ=M�J=C?�&�=��X>�pνC��-Z?kg2=�s5��=�9A>A6$�{��H���H�L�I>B�>[�>�:>].h�:��>u9H=�v=Wq?�?�ݺ>q?޿�a���ɾjx>���><�m>�w>vCA?s=�>��[�����>�M5>���>) �>��;SP��l�>Ӧ<�Kb�=�$>ɢ�I�����=>����k�*>�H?9N ?<��=�c���0�N�9��[T����>j���c���I� �>�ɽt�=�Q�<d��>�����@(�=�Y0,?c���5��� ��k�>g���?m��:ʗ��"8�=���@�����9�>�����^.�H������>S�9>z����>ǧ��/XW��l�}'9�r�>>7��>9�<~<�;.k�����Э>�@�R.þd� �O�J����`�>�'Ͼ��_mx>�Խ��g=�湾̎�=}(��k�M��#�a�	�ۿX?M��K���D��e���A>"��2D=�?�-�>,����+Ӡ�thV?i9�>NW|>��u� �#�Fk�w�.��!�>�0�<wH �y?��=��l>�N�;�>��>����R��=�R�>[b;>��y�̰�<:�Z� >B���>�f"?e&���X{=����)>h��������> ��=�*:� �K���'>�S
>�T�>#Et�`2̽�6���.�m��<�e�>�>�:3�+���#��Ň>YoĽ��>K+�>�h>-�o>��<<���=G_��Y_����Q���r?b>�>&��Q�,��"��$*�t#H�bh �d�y�7���*�?-ž���ּ۽!-��|�����p? J\>\�/?U�Y����=;?���<����.���7>Zt�諬>Dؘ�D2�>i��&�F���]>�>&?*>$nP��E����*�[�>w(��v#����>T۾T2�>��C<b��>f���փ�<�v/>��K�����,�?��?(��3����<u��|汾�W?��(��=6���c�>�R�A\����=|�=ֽ����p[?+�>��L�G:��^�=������q��>��>�Cྱ����䄽 t缵0P�>�C>�&E?#���V���J���-�<�����ܲ���A>YC��]���{��Q޽d�]?�8>��w?!�Q`?��c��������>�jн� �oђ�@�d�z6�[���䢵>� ���_����,�ȼ�e�>�f<<sN?�b�>Ӳ��Q���ľ�J��	��>��3�����\>�灾��p> ����=�"?N>�>��x>/š�o82����>��=�ۆ��#s�����3H�>U6�=�좾�.?`�>��=Y�N����>}\.?�s>?C���\뾛�<p]�:��>���l�>(�u��ug�,��>Nɽ�A8?g�r?>�>B��>b�n=����ܜ�>�ζ>���>�$>?d��;��$>=����-��s��>�s�=�>�ʾ8�Ͼ-�	<�|���U�k/�>��	>���<��f�ʾxO>nk �|@���?z�=�6�M����S?F�?,Y?�2>�H��.���|�>m�P>�q>d������>�X������W=;��>QѦ>��S���b�W6E��'��W�}>P�>h�پ��>>n;őL>�䷾� ?a��>�Ɯ>�,=&-1�="�je��|B��b헾�]�#CW�ض)�����	@���z>^�{=�������R��(�]���P�#?�j��P��= ��S��=��'�w��>(�em=7x&��=��ٽ������S>� �=B�=���>� �>�E�h'���7$���<�o޾�#?%۾8I�<�b�
�;�Q�d�>��
�/��@���0u��̫������T�T=H�{���c>>1�־%��3˽�;��n��Q�a>wP
�	,>|��=q4��ލ >�t�>�Ŝ��1.��e���x�>��=������S��L�x$�ZF��#׼c��`@2?ޯ�>�R(�\�>��<�N>���>mJ�=B�?�),�����=��*q?�˚=J�ܾ�;ҺA�>����]�Zr�=�/v�����0�:�L/��FN?V��lľ����zI��Y��2@���>���=�W:>ڂE>؎>\ >躾��V?�yk>z[	�0�9��1�>u�r=M��a�`>P+2>)��>��=���=0��> N�=�Rj>����y�<$�?{����'=U}>� �>�X�������d�a����x>��=���>n�1!�=�d[>�z��v���=���>�~>Z���$������|/���zr>��$?��>�=��d�>�AO�>��M��$�?i�
?�S��o��a>�	|�b��%�o�F7��䊜>�(�>��B�.9����&�>]����۾2 ?Rb>I>�9y��,?X�e?wq%?�����}�>�ᾴK?[k���z�x͎=����Zhc��s�>�D>�be ��E�E2�3J��؀>�h�>p">3�����r>s�ʼ4�X=��Ҿ�?\<�=)m���ý�I�=K�<p2���L�>j��=�� ?=c|�����X?�%>��l�0͜��ĥ=;�\���%��>��g���g?>�_�=�5?xv>/�&>�Ta=�g?�D�=~��=4�=L�=�]-�>��>J&�>������=�8u�>Zn?�t�>�����[�N��>�\�=ŜD��p�>#ٽI&>_S����?x��>l)�>�gѾ{�ܞ˾�I����^ݾ�;�>l��>��>Uo3��5�<oR�=Ł>w���9?�5?ຌ>��ic�w���>v㙾27����z>�/a�D3(<�?/>w3>ZW����>D�??(	?��<����"t=��ξ1E�������>w{�=`��d����ľ���>PR{��d�Q�>	=�2d�GШ�΁?�b"?#�?	s���6�=:#�>Ȁ�G��/�R��)�=��Qsɾ��>�Y����V�����>����r���|f=R���̽c�)>k�C>�><4@��R(>z�?�	��{B���>v��>F*w����[���G�d������23�!ɧ�n����>�]�#���;F���=��*�$c��#9V��b@�>F�������=ܾ?s���S ����=��i��t��H�=;v���*{�Jǽ>��c? �>!�$>�!��vp�;����+>����6�>�?%>鲾���Ⱦi
?�R�>��>��H���%��d-<Q<�q!9=��h�/���>l�V>?+��y`>��>�>���<��=>�:�>$al�C��<]����><
a��j��C>B�>f��>�����=�Q8?��1��������=8�>��6�_���-����9��;�ZJ�>�El�
ZG��_|��վ���=�=<��<��{��ʺ>Ѥ�r�?I�<>1��>��Ӽ.�ǽ���'�>�};�����`>!>Ľ�p��By��?�H�V1q�Q� ���>�|�;�N�>h��>��$>��>xf">AB�>k�?`֭>���<-�Z>��)�<ϡ>�!�Z���6��>�T������ޞ��/)?�g�>Z�o���>�:!?{�*>R-K=��`;Z�>E�վ����b�9���>�z\�1�����Q>�|;>"q�>��T��,M>>�>@��`�k��Iý�>
+=�?'��u�%�����&��c뾐@оe ?C��q|C=aZ=�)���Y�=|���_���>]?&��;2{��7�륺�<�]>T�;�=>�OO�� �>��>��r>�?���=x�>�qz�9>�d�>�I½b��>'�/>�����^?�6���:�G��=^Ӥ>ɱ�<�4�߿��0�U凾F�;��&���>��P?�E�>&.>���=�O}�T���g�>j�>ev�>�7y=�Ӊ����>,֬=Bؽ>o�<�	�>��]?�������=��>�v>�>���P�>d���D>��ھ2��>3�?%�=��=w��=7���6�P����>8�j�*A�>>!�>b�-�Q?�f|�>��뽝��_aܾ2w��戾�e쾥�����?�L?��>>\P�	��Hh>�G�>�p־�Q�>/�T�_(���fr>�s�=�8�>{~�>PT,���?��ٵ?[�3>K�>��߽�5�=!R��촯>���%��=&��D;��+��rt=�����Ӏ?���c�=sϏ�;�1�u��>K��^{��ٗ��k�t��>n?a����þ��>~p�=W��h�>�����d�e��Ǳ�> ~�A$޾����`>8^ɾ���X�?
�?�cݼ�М�"� ��W�����>X�?�阾䜄�Ƅw>�\1�l���H��6�>���74?�8���<v����'�M�;��l�+C!�ڣ޾IϜ>8��> �i�\��n;���H<K� ���U���z?&~�*�(�7�F�Sm=G���ú>��ﾟ�T;��S;@y�>`�N��a��=7��\�>�r
>��2?(�>3/�#N�>�L����_��`�@�ϔ>��{� �1�u(��ދ>ik=	�	�k�������Q�~ނ�fdѽ�-��kC>B�>��ܾ~4�a�=�⤻qWƾ�S����M��1>�dܾ��,.�>�/?p���ؕ�yT�>��@�6��u��>�`>�����`;�����-�y��٦-�)��%
p<Ԏ	�2}
�~���k>ʾ�==7�=f|�a�O>8νm%�>$+u�p�����>iS���z����>�l�>?��>S�=٨z?�a½*oྭ�پk���Fѽ�J����G�
>SX>�>��Խ�M?�F򾨩�;E�ѩ��X��L�|>碔��饼8�P���B>�j�>4��?[���/D%>�ֹ��hs>�(Ͻ0����)O�A��G���k4�>��=q�����ͽ9^>J��>A�?Ee����>|"�>t����>3ո����>_>���u�ȼ�?8
��]��H�����
=Ho����ƾN5�>m�7�P�>nz�>��?>ȣ>YU?��>L`�=�
c?�gA����,#��~��>1܊? �>�>����M?
H�>l�=c�U?��?(���q�ʾ�d>��=g�>tV>������>�=��I���?w��=�?#=��>��7��|<��Y>�=Evm�q3��³�� >��L��i�7� �� !>�:p��KK4�b���oCE=r�>��ʽ�B̾
��=2z>Cz�=nAݾUӽo��>u(�="᩾p��>��^�URG?D�?� �7i;>�	?�u���>j��>rH?�%��qo�>X�>��O��m`��=��-��YBh=k�ؽ�����1��2?�=���=��@�ʷ�>���>��?)�)�U��> �=����7�V?>�_��ɾ�p���׾�(��Q��>�So�΢I>sC����?����j;�=B~
��i�����q��>>
`��>C�� ���P2<�ё>v�#?���>a�ּz>�)$?q�>!w�>�8c?I˖�8�~?~-?�T7>+BF?T�%?F�|>c|�>�t�>�]/?H�m?%�L?�[v>�>���>�o?{���f�A��a��]��;'�A>a!�("�(ď��$>�B��m��t��z��u��"����0���4�����<��Ǚ=��Ӿ1a¾PC��/m�<� Z��<?���^#��V;��>4##�q-��a����ۼ�8����a>+�=�=�~��m?2 t>�_�>��>��o>�@�>]w?t���A>�6~�P�Q=P��>�WZ>)D	=A^�= ��i��{O>T锾X̾o��;�߾074�L�*>]�?���>v*>n��>�C��ț��~>Q�A�Z}�>T^�<�?��j>���>b�?G�>W���)�&>�\&�a���վ��=� > T�>0.�"P>��;u�\>��Q�)y�7�$��g�>�څ�����#z��m>�` >C�о�?�>�(�d�1�湠���p��ʚ>#J>��&����~�(�uu�-�
>��j��T�>C�E>\��>KF�>g"��%��xo�>����l����io��9>����#�j�M��F�h,�=��>������b�Y>����=�g>�#|��1�V>0�2>ž��@�>+6h>K4��B-��]������>�_o��(��l�D��4C>�읾j�6�'�#��d�=A^�<p�<>��9��
V>|��J����ݾ�|U>)yS>�e���>}%�>Y��7 �þy�?��/!�����4뽪N�>���?,
��`�=+#�>{���<7�>2�f=�� �w���粆>2�>�Nٽ}�8�A��>��?'���#w�>Xd>va�	�<�������`J?�̼��,����=��^>���fA˽���>����}ؾ��M?T���Y���V�?�Y�O1�>a��}$?U�k>ʹ?�Ҏ���?/~����?�����<�V�U�?���>Kk
<�������>Ww*�f�� �>{t�?���>��>��=�e�?A�޽��#����	>#]�����0���<�k�.A@��aɾ���=�֐>uQ,>-&I�ŵ�=DD�u韾:u���lC>9s�=�3?k>�񑚽���=\Z�=�9>��t�sf>��>� ^��ˏ=\��>�B�>�?Z�����&��=�彩�>�_C=%=�O���g���k�>�?N�4y� �C��q;)LH�a�;>i	���T�=g�>�,{�Wg����Є��;�>�|�<Z;��ǂ�:�ɽD������>�Σ?��y��6�9����5@?!x��,�?���.r<�O^>8x>?*�2>.�>z��hA�?��=�l#?�\��YE�>R�C�c��=ب���g>�b���E����?�p�>�%Ȼ�̎�e���D�=?��r>ul�>l�?�Ӈ=�&?r_?�~�>(#d>禅=�[I?�Bz?��H?Ύ�>�w�>4v�>ρE?�r��~��>��?1,A>	�%����>��>:!�>�j>�c�>_��>�.�>����a>l�
?��
>[���4���]�p%�>�GԾ�~M�������>�$�0�^��sA�z����9��=A��q�j<2�?���*���T�6u���-�Q��=6�a>D"5�sCV�<]D���$>2��>�
�!b�>Aa�>|U��_(>��=���>ac�� �����=$7�>I>�@>f�>���>٢>�о��0�.?�>���z>1��>q�>�9��?�;�Ե��k>1'�>Ԝ����	�@�>btU?V�A>�튽�����?R+<%Z�����H�Q 8��$7���%���W�L�h�1��J����:�mӾ�4��uEϾ#�.� :Q>v�sʾ|�>��>T_�����&�5>Բ��3
�g�4���8�� o��Ke���ֽ���>z)��cO�=	h��Z�=�d��	)3?5߄��2>82>�;�?�����=���(��?hZ4�^��H���s=�Vg�ߐM���x�!�B=����ҍ�۷��	x۽��=?Bv���Or�aCξ���>
ч��j�C`�EӴ>�ž;w����}������E����о� �>�3�&�K���=� ??��>��E?a�>�-�>K�k��-�>GU>>\8�>���Yr�^>��`?����_�>�V���?9��!�0=���=��I��/˾�Q���x����³�<�6��Kk���ɽ��A�)�{�F<!�)9?}��>���d5L>����	�!k>�P�>{�?�?ڽ��K�w�f?�)&>�5�>�|F:c	7?��2n�>.�׾�����d���!?|�Խ��ܻ:3j��>���>� ���¯��*��n)�OL>��>l�����zx/>O2�>�CɽX�l=�+������o����SZ�5/|>qV1�ڑN�����J��=�p=��&>
f ?�%ǽ=|1�%�>�>��5=��U�q#>��>�S>�tw>�㑾(�?����/,>S;=:b>����L~C>E�>�㽮��$;f=��B>R	E�Z��3���Y��]5վ���>p�ǽG��=���>�ې>|Sw�P�=��S=�3>pf3��)(���`>�>�4=�Ö�I��>A��=�</Y>�?7Z���=sw�=(n�>�m���<A�e��8?�qZ=8��=�ܽ�2�>��>�,0=��u>i_O?�,>����>1��>g묽9�"�>���|�?�T=����u���?Ny�ˎ���>j��/T��ǎ�>���=�!]��Wt��,,>P¾>�>��Fc��G����:�= u��t�=N������K��(�>'hȾ����y�����>lD��m�2%L���?z�>�x>%�>��>j�o�]8(�$[�L3~>6f����澁����w�>���>�4i���_��?0�=��>���>;�0���b=}�n>x�쾸S��wQ<>P�����&H7��ǎ>�*`�a����\�=;{���C>��޾ϛ>�~��V����m<IE4>��C�^�6!�Q�?�+ӽ��^��#�u��>�
>�	=��=�*�f�>_(4>5��=�����=���>d�=7Y�F(E�ȝ!>CO1�G	¾�^����cŔ��=?t�P���=�k�>0y�>� ͽ�+���=r �>��b�DV�O�J>7�=>�0=���<?�>5Z�>T�>�!>)
�>q��<`SV�+�h<b�=�In�Kzy=�ҧ���=�].>�ἅ >} k>���>$%3�"Z7���W>��>V9x�v�s�L�Q�:�>�n�=r�ҾW>R�>�$�>bW>E�> �2=I��B>Ֆ��t?��B�#>���5�M��w��b�'I���b��ql��Y���2�-<P�޾��|�V�y>�{S>�+7>��C�i4���p
?�R�>�N��j1���!>A�(>�+�T�<Gt�$wE=+0�����=�;w=^}>��'>5�l>��ɽ(f?{�T�q�V�"�>B�<��=m�>H�>����/%��L(:[
ؽ;�!�q]O�5�R>�'>x3��>��>�{>$���N�I�)Qr�O��<�z�����=:k��|�e>��W?}�μ���0|��ţ�>-2���>�D\����>��W>+��>���=���>�I��MݽN"�W,�IOk�K�	��z=2�����7���>��M>�{2�>�i��?����>�=���l����= y���~�,�_�#�>jB5>�b��ؖ��N02<Qľ>�祾d��ٓC��z����ͦ>*�`;+�=w@�>��>��x�������=a�v>m��=�����u<>���>i2�>��>���>�f㾽�þ��׾����
;�o ���1S=?ȽH ����=D^S>�6�=�L����>jj[��6�=y����n>�ؼ���@;����=f�*>|\>T���ۂ�<��>\>?�b�-],=)牽��.��~����g>�
u�j{���|��G�������=hxV>��=���>�(�=z�T=��:>�ϯ�۔	?��,>�~e>�I�>G��>L+=��X>�x=���>���>s���̕��>I�7>M��=����^��q�o�=��w<&o���ھ��<�I>�!�=������>~�?��ռ��K�*�x�M<� ���>������<슏>�+�>1Β�Hǽ��н���>����:�=�>�t>��L�0aY>0�=ba>��B��#ྸ	>@�%>�>�����>��>�>{оn����]S=RD��&���fu�H��ac���1��x>����ӿ�S��="�O>Oh�>��ž"C½SF�;��!>�T��o�&�>����9>�x�>��xU)�(���G?�L=?3M��5B�$�8�N5y�pL>�2'�Hm>�������j����Ⱦ�:�)�=������:C�>�[$>G2>�:G��.V=��a<�.�>փ꾗����s"���?��S������>섇�k��?>L�M>�m�>c���t�-��<��o>�!�����>���v��<�Q=�Cp�=q�W���x>�a1���+�!��=ɏ������F�&=9r\�?��=Z�nC�>�H!�2��0�)���=> _;�	޾�����>�0Q>��ݽ'2�ݬ6?�=�]?k�ؽH1޽�p=<�A�=W5��Zm���=3��H�Z%۾DN���ٽpS��ܘ��ž6d�2�_�?�5>RY�>�1?��0>�9\�_�� ?�>绸��Z��[��>�G<�1�=�`M��?!��>� r����=�,�>��>�n�<(k����#=��M>"Z���J���>��>B���W><�!N>���I�/>�[�>��>Q1�����>�e=�Xb>P\��؈�{gH<��	=%	��N/ ��dW����1�~>A>_馽⥾5�t=9�'>uT�<C/���E�=�Eq<k#>��i���z=���,��=�ར�f���>� �=�T>�3��F�=��k>���>�c��7��|f^>p&>>��������վ���=����}=��=r��*��*�>�#R�>�F�˹��t�WV%>@0�CqF�;�=��پ�k�>�S=="��"]?]=>�#f�>�#�Df�>O>�����ȥ�U]�>V�=9&)>S�ͽϟ�>j�>g�1���#=E� >�¾>�k��W��[la>�w�>�=�gS�EA�>E�>q��>�O
>���>H�z>l�>jrS��߃>��)��˾���>�$���@>%dP��!�>���>%��-}����=�LV><%K=L�E<QDb��Z>M�>��1=�/1�	U�<���>Vc���#��6�=�Z���>�Z�O�#>�9�=;�L>?�>� �g�N�bS~>q�?�oʾj�t�����?���m�a����}?����¥�=��^=(�=�"����v��>�q��ؽ��P5�<$?>r ��J���A
��&>������F2>�Ъ���G�6�˾���`N(>��<"����<[>��?9��6��` Խ�5Լ��H�}ɾ#���I�=�u��aǪ�|T�>��>$���w���S�=/<�>��x��!F�Р ���=�����G�>AK��K�=�G>٣�>���:%���ab<C�|>�C:��%���<���=+=L9�p=�">X^��0N>�F½v7*�-���X.>�(p��r�P=m=���;�?��v%��-P��T�>,յ�]^�����=�(���"��
w����=`��<�ӭ���]�z9>��>�<�>}��S���>���vT��8'�=F��<r :>����ʜ<R��>��#>�"�F��Nk�>R��=v�о�݅��B����mG�>�B��a=��J>��>�o4�E��֓��黛>-t �j:�9(O;�;�=B�>��p=�C3>K�>��]�p=�A.> !�>Dǻ�/�sw���A=mX�;/$�[��<j��=�=<W~��ۇ=t'� Z�=��,��n>�d�������v|=r(?�{�����M�r����>VO3����;5���.?GU�>W���֟��Y�X��>�	��pá�?���	?!��=�a �������>�>�%=�ќ>�`�>�|�=}v=+?��>������U=|�����=��4>w�����>���>=%>>>Jy�>�t�>���=�]	�I�ݽ;�0=ζJ=E��N����?SB�=��+�'�^�56�>r�m�-��>�L���[ >-r���zZ�Fӧ��C�=�c=� v����]¾>�H�<�}b����C��>���=ڲ	?�^%�'���w�
��i,b���׽���=�����F���>R^�<+��=�j
�S%ƽ�gg>!�>F�ҽ�O�=��}<��]>�ˣ=��ѽ8#Q�h͍>b��>�Ǿ֣��٪=� �>�`վlT�0����ڧ>ޔ:?��%������3?�E�<a$0�3p�?��cӽ�h�*���Ld��ƥ=ܘ�=["q����� ?�?��1�*���l?��>�H���,�>�A?���=��m��?G?��>���=��=�0V?��>=Ɲ>�J�>�K?6%?i7�����=Y%~><��>��ﾴ+4���=��>O�qݥ���L�<<��?��>W����*?b�����&��~=A��>קJ��
��~>�:�;�x>��>��I>^?y�k����>=e?�?%B���O��~>�?��Y�]<��l>��?j^�K4������M>��?��?tw�=p�g?�Vy��h��"�>��%?	I����(�sT.>=��;�P�w��>�z�=�:�=Oi��^��=v ?6�¼qi|��c>�y�>kw>8W��a�<���>���>���<胾�		���V���y�>m������F�Ҿ�W+?�x��̾Px��v=>�$�>�b½%� �&�+=T%�?�? 
�>�-[?x>h�'�o����?g>������+!��t�>���>c��C����I>tVE?	�=H��ۡ�H�j�ܵ�>�`!�����g�#?�J�>�Im�đ>ŤؼXmξC�>i!:���3w"�Z˿���1>>2�}�r��M�{F�>L�վ��K�γ��	p�>��=��#�A�~����>Qps?�AU>7վO�;��2��j?�E�G'�L�=V�">t����	��ꂣ���H>&>�����e貾��9��i]�
^�>�x��pʾ�C�>����3P"���w�O�> ڪ��`��u��"&=Xu�>��>=a=�I�=�xJ?3:�>[��=#@u?=�#�s�E��`s>���>Ӿz�&ڽ�38�����^.>���=��v��j���6�>[i>������O>VЂ>��>4�Y�a�%>z��=X�{=���析��_�>Z��>q֙>:u?�3>���?�ng>�>���>�G����+��Y��Ѽ�=� �}��*����K��ӣ�%G?�����=2S7?�n?q���0 �>�3=E�?[W6�����%��>yt�>��B�P� �&*�04�>͘���P'�p�>G@�=����I�*?#c��\�=ַ����r�[5'=�>
>�<������=sY0?��>����->��?���T>!�?X�>5�v�N��>8>O災�k\�PΊ=z@1��`ev�S��>��>ww���7?yy���'��r��>�*q?�S�����7B�>2i? ��<��"�-E?�&�?�:>�t)��E��t��� �=-4�>�s?��¾j��;�mg>�n�>����:%�`����>�D��K�Q�AI��hSa?��׾��"�t��>ְ>�إ��<�<�l^��'�>�_��sJ��U-�=H
��!?����<�V�=�稾��<H�>�p�=�����)�č�>� S>�.��de9�r>o)�><t?�8!?{X4�e�Z���Ta����>�Hu>h�?��½nr�>�o>#+A?�r�;a�R>
�1?2��;(F�1?��z?)*|��˪��j�>�P>���?}-2��+�'>	vQ?KݾW�^�b⿾�u�>��G��>
�� ����v|?�$C?;_�����>h�+>r�>h�>��m>��>��>�� ?�d�<�X>l?l��?�~?��=H�=('�=���>�UҾI5>U�S=N�>Ѭ�>����y>~�6���!���%?q�?��ѾC�O��<?Ą�>�u?���=��=�=�>�y?����m�C�P	>p�?��T�د�c��>����c1�x�¾��T�hzu��s�q[�������(�>*�	?],>�!>��.�=�?�j�����>�)?��<�Y#�*ہ>Ud>�Q1��R�n;�>*�>gJ0����D��Eﾝ�5��y���G�>U/?��e�����>G�>�<ؽS���Kgս|��tJ�Q�>��>K(Ҿ �U��_�>4����2�n%�>�>�S#���R���H��>}D^��cG�	�H>&��>l�
��	T����Y4�|F2?l�,>0�
�󉕾�:9>���>æ0�w�*>`o4>J:�>}�6>�ߗ=���Wﾜ��=�eH�{��=��O?h�	�٥��Ò>hV�=z���Y(>��4��߾\Kh�
�1=�!g?S�>�Zn>PX�=��//��)3��Gt���>�\ξ�@=�)����_>&US�k]Q��N��4?��>J���k%�U&�>�cؾ�R�=v�7�A&?���>ھ�~�Y�/>�&!?�����^��]Hk�8�>�y?�%��s�=��w��[���D���=,�F�7>�C�qD�k�w�n.оG�ٽ}q�>!�+>�N>� ?g�޾}�����33�>a������D/,��R>/`�=T�սVý�tw=�>�ɽ�C����>��|�q����4����>V]�����n 罨��C�>��>��7>�&�=(kc>x�g>e:?9 �?;B����=�z�>�0 ?�$s�A��ʦ���%?:���U�J�n��*>jL+>U��>��?R����? 3?/�flB��HK�Y�>{݇����a2=M�ϯ���}��z���"�>8�?0�k�у�8n�>5�V>	8�?ʚQ��Ko��fZ>�!?����.��aO=ڌ>(���j?��P?bbe������ݽp�����<l�H���=��S� ?Q6�=����a�%`?d��=����%2�'&#?(����1Ⱦ�82���>��齘y��W�F�	PQ�VX�=�_>]�O>��=>�=f�
=�p��V���:?��$��Ka��6~�>��9=�H-��$ �A}z>���>�aK?���>��9?��Ƚ^(�>ɷL? �O�ߨ��9�>E }����>��<>-�>�����	?"j�>��"���ؾ����8x>r�>?�n��A�}<b��>ԯ�=C�:�RK�>�פ>z�9������ 	=�d�<�CI�	v�9�N����>
�(?H��>X�������3>�8y?;� �y�2�[>|W#?��&���������>��}>�l�>ҧ->�W�>;�KW�>��>�l�>������%>�cO>�>�xY�χ>Yx�����;���?�?A��>N���:'H��9?�c�>3�>o�d=>�G>�"�>5}��c�������=��� qp�dI%>�{߾�tT�.�>yjH?��M�6�=�+�=O:D>���>�i�n�;*�8>_=�� ???�P��:��U%?�5����/پ�x���~��NQ��eξ%+Ⱦ\]^>���>tB����g�10V��x��Pf��A/�$�(>2?*��󽫏6>6�><Ǿ'�?��,�%���˽Xp�=Cݙ���6�"�.��-E�:�>O�>���>l9g�Y�5>�!�>	'�>�Ay<�_d�u��I�>��o>��}�Y��> )>m)|>h�`�Q����>x�x?�+�4Fʽ㣝>��T>�_L�ŝ�Vy-�،����$?J8�=$��$�>m]���%���ھ�U���M����R��R���ӾNz?��g>A��<��!�<�<?�U���;�"f?O	��V�<󭾲3����ߴ��}�����I��><ŏ>~)�ؾ���>��S?����>~?Y���1��(�<��?H���1AM�� ?>˿>�k��8,>D�?�<E?�6?�t��\���Z<���>��
�B���*?��ʤ>Xb�=��ܾ�2<��o�>��[?Jmj>��f<S~?�! >�ݜ>�[?���,᪽�/�>���>l]?�Y>��>
it�IM?¢p>�_;��v	���?�w*>+B�E�z>���>���O�4>�$=�J=�><{>hX����W�lw�>�t>}� ����i�>�Qb�4�e��sg>=��>�	��x-�L9v�{p�=9�=�[�>�۾�A�=���>C9?��y>���T����뾰����!�>���>��о��v��(*>�o�>+�>�LL����>
r�>mf�>ӳ�\"�>� R�� %?� D>�A'����SL?P��>Z���Z����>�׎�������.�`n��L�|�z?���>|� �y�>?N�>��M�Q����>��6�;T�>�X��2t�=�L��d)-��Xj��9:�_^;?��r?{A��X�>��v?C!?�1?��F?���?O��>��>�! ?�&?�q�?��>�� ?�_�ʝ�=�JԼ��_>0AR?3�Z?}<�>��I?œ?ֻ?�\?� ���u?�ÿ��ſ���>^E�?�q�?񕟿dP&?Bȿ]�r��j/�RD.>6�ʾ�xZ�Ls���?�ID?^]���Y���]f����=�r"?��>9��=�4C����?}��W�(?����5����D�>OØ?��>I�þ:R0���$>o�C??@1�?�;?Y�?��qԾ�`P�ۧ?b�UO�>���_�=_>�e�>̾�@?1�}>$��=�a?O�S��P>ğ�>7�?��>C�4���N�r�=�=@�z�q��x��*Ž"�������p�_�.>L�ž�_�?�ㇿ��H�9���rh��d p�@����>s֣��~ ?S��<�����h?A?�t>rI��)��͏��N!�t�Ҿڣ?{����W ����=R��#�r?\��?ʃ�� ��r�տnk=��㘾[6���Ro��g�ak��fN=�;�l��>OҼd�@������Ȝ��e�Ӽ??:I>��\��C�>)�Z>��V����͆��?N���>��C�"m���f?~�|���ž���>��>�����>։���v�0L?�7]�j?�>숖=��<�2;?k��r�Q����t�)�.���(?��.>!���ٯK?^fν��%�� ��؟�]JR>�Ŀ;jYɿDf�>8o?����G%D�B�>7��?�1?�U��6w?Dh������&�>���=���=��K�}<��5��>���=�&r�9��47]>�%ڽB�P���Z��N?y�8��!)�@���m>�Α<�&��r���n?ԏO?���?|�	�bst?��v?7�&?���?Ͱ;4����y��[��G��'�����U?�`�p=���P��d�ޟ�M�=�_��\?Z��?��=��A��?��?p��>R�h�=�#?aD?�jҽJ��3D?��:>��=��<���7��ΝƼ�"?>%�=�hf�̚�>�k���=��??E���7?��Y�В0>�3��=�?R���"�>�Bn��cp�e���H>h����i�?4G]>O�D>� =�{����=�E'?���=G�R;�BH?�_5;E(>���? ~%�"Q��ո�>-�⾼�l>N�����?�D	>y�>W��l$��BF?R{�>%�?<���2���
�>9(�?�?@�/�8=�v��:?�EU�'��b�g��tɾWI�=7:��e��D$?��־���=xiG?m��<�<�M5R>V��x"?�Ƥ�������vC?���=�S�=h���Y,����/.���v�w=�����>s̐�y�9��|3���C?� ?ˍ�?�I�>�$�>�ȇ��BϾOy�?���WV��=!g?�em�3D����9P�<rMH����(e�>ik?��?6sd>�|u�fɾRՂ?|ܾ#!�=_�?w�r>eM�ndY>�0>�f4?2���"^d�7�?c�N=Dŕ�V��?�n@�->���=p�>�?��<?�u�_� ���-�q
���>��s���N?�L�?������.?��>�s�>�#� ��@^?~9�=��=��8��:�=��*��(?��������u?X�ƾ`'��Ц>驾?w���˂>P
!?I�"=ʞ���о0�>Sa�>�9�>3�)>�>],?!ۺ����>�">�H�w?�D�>wI޾[�y��vľ��E��� ��'���[ּp:�[[A��-O����;5P���þ��H�V
�G��?DC+���?��XP���	�-}��1Ҿ)Ġ��Jſ���r�p�;埿���c۾��3���8?�\??s��?J�����&>�0�=Wʭ?�C���J>]��>\��?m�_�%�?�A> f�-�t�`M����[΢�\rc��4k�K'�V9��q��/͊=ٸ�pˬ�Y��>uc<�V꾡�Ľ	:>?��=s �����?�)�%�?�Y񾽒^?Z$۾�9�P=�>��U>j��><�!����2�C�<.����>lTq?���>���I?=Z�횵�AW���H�� �,��=��S�eݱ��3X�6aս�&��=徭l�>}e;�MS?fz��mӾ�Vc�[����6��e��I�=,ss�*�����Կ�=��\���?�տ﷿PQ>ޅ�>�O����0,��9)Z>�}��:�g��A=��t��ZX����>�@���u|�y�4�H��<��>HN�����?>)��쑿ꡃ?�s�=�R��u�?���>U)�!�?��Ⱦ���3����>B>���,.a�z������?(+�>��(>��	=�)i<&�V?�?C����1?wK�&�j�.��\w��y�e�;�������f��<�J�P슿 7��;�?�?0���7:?��Խ�?W��<�v�>�0ȾW�}?H>N?L=��
��o+ƿ�䁿V�>קm�~�i=C�=>'�]��:���k�?�W�>�/�N|�>3O�� �m���>����s;�5?o�������V�?��?a�j>R*���І?��B?*�=��� J?���?��?u��QF�?K��?��?�>{g�>�w��i��Y�>��>��;�(*N>���?o�?As�>O?>�>��=�l>�0Y�1`q�����k�*��3��23?�ֿ=���a�޿-?R���ވ�DvD�s��>��?6c�>��ƾ`y�?�㧾���=��->(���)���e���d�z�r>���Y��=��.�{�2>�~�?:�>=YJp?0�?lQ��{>� '>૪>Վ��~R;�R[?�\.?�?o��u���A������W�OO?~�>= �/孾B��>����Z(>���>M#��B
�>a�>��>���>���'T��%�˾�.?R8���^=�q?Ϯ�?3ϒ���<��?���>��6>血����>�o�?�7e?ٗɻ�6�>"�w>D(�>gfX���H?��>VY��qޘ?�Q? �?�����ۿsv7?�%J?��>�Շ��
2�%��V�v�@/�~w�>qpg?�켾r^>^Q�>�7>ގ��M�z��>��9?�5>B��>գ�>a�?��=Kw�����>9	"?!��a����J�>L�?�/�<�.�ҭ?x:?�5�� j�=��Z>��?�aC����>��>�@ ���@>�jK�;ri�%$f�E�?]>s=��ھ����`J�����>���kH��ò���>�~��x��������@�8?���>��I�Z�>��'���?]ƾ�9-���>`���v��(̓>12���o�?b7����˾�Q�<^��>hۅ�S���� Y>���?r=�a��>9�>A?�{�=4䢾�ʈ?k}K�a<?~�"��jO?0��>��'?������T?�N�>"?��(�؈�=d+>�6�>�,>>�ͅ��r��B��>@Ri�%��1�G>��L?���>+@Ⱦ~�ھ�a�&`��о��&��1j=o�? (�<�#
��C�<���>R��,��O�=WO�i�!>Ⱦ��<�<��8O��Ow�%��v߾��?3�&��D>�4�>A�%>�?�=��d��X�=λ>	?k�_?�<��5�>�}G�t��>
��<���7����=��>��ھ~Θ�Z<F�3�B>}9��r���70�>�����m*���N���	>�k
?~��>�&�&�Q?8�8>ȋv��I��|>SM_?�2Ѿ��߾�7I��IU?hɿ#Z��$?@ט?�
{?�d��_?m1�?��t����㽗?�	�?����/|������I=��>��,��!Ծj$o?�������o�S�>D��6�B�$R�>IԾ99��F��g�C�����=cF�� ���i=� H>ݫ�6Da�����d��Q�>��$����?����J$�r:?�ju���??�?o�W>��Ͼ�c=��=��x2˾*��?k�!�� }?�8>��n�?��q>2O�>�3�����iؾ
p>z%>t�?�<����>�,?\�输�>���3(����S�ʕ�D�U��A8�L��Ggl�l�<�Z]C<��>�+�=��>�"���M=��<�e�?��S?v>p�=��>�#T?�{?-wA?Zx�>r�C?)7�>�A{�M���-Q>�2?�tY?4$�W`�x��=�W�45��D>����i������=>"?�?�Z|�?��?�y/>�^��e>�蟾C(�%�I�E��G��u�;�Um�xl?I��=���>�i��R�>c�ھ%|�>�Gb?�D?��}���Z��TҾ�=I�����$�˽�~���lt>14+?ݝ�=�?'�(?�s�>����	?\?=@9��[�=ѓ~�-��=�}>��M�78?��	?Nlk�-_߼&Ծ�~�<^��>y40?���wv��G�>듢>yTo�����dѾ�´<e־�D�I�j�@��a��=�能��h�%h���ǽn�?@���p�#ZW���h?�<�>��=�}�>!t��>t꽶�m�n�x?s���:dֽ�+�,�j>��g��>��߽�"��Kmv��\���e�����>(홺.Mu>}V��(���r���>�.���)�+�4=����Y�>�������w!>���=d@��|<�N,�ځQ���>`� �z�|���=�ՋC?+��DQ>�a)�q,?yW�o��a~'=mx�>��?>�#T�]̾��S�"Á>��>��>����4��&F����=/'�������{��,0�А�=���>buʾt��?�?���=�'m�$?硽��a����~9��z��>���>
�.��.?��x>��e?|=a>ə`?x ?�jܾY�Y=8S��p�V��<^���-� ����K����[�3?�AY�]f�=�_�̂�?5<+���=$��� 
�>�\>�9ݾ���>o?�ƣ>V��>I��=���>������>��e�[�K?=�
>(����>W��=�w���>'۽k�8�.ɾ�J���|s�ɋ�d{;>�t ��tZ�YS!�N4=�/�>�ʶ>P����'I�gQ�ֳ!>ks�����r�>�٪���>�ݢ�G&:��Ł�� ���=�	F>�'?
vf�wR��O3����>�ER�;eվzN�>R~���>���=q�0?��G�U��=^�F�h?������>�2/?�#� M�>t��岕>
�X������-�ξ"6\?���i��=%�7���>W�?��S����==� �<$�{>y-��］װ1��!��GW9>�s#�� 6>�G��W>?C�l�T>�=��>M�j>��,���=Op{�"6���O�<�V>�2���S�;X��'�9�?|�>���/�>�"��ꦾ��<�䀼��վY��=A˾���"$��*=c?��h����90��>'��>�a��I�@�]>�&�> ��>�݈>L��>M����e����(Q������Ǜ�Ҳ��>��d?�0?��a>��?Fi�>���>��>M]��q}?��ӽEC�>e*[=��$�h(+?ߠ}=<,g>򨋾�J�=��6��|?��������>^S�=���=}�����>ljԾ��\�|�=#����?F��>8�)<�z>e@�>HS~>�'>A7�?�XF>�nB>Ȋy>ϰC?�kּ��<?�>-�v>�D.?��a��Ҿ�`K�/uB�'>'���q��m�V�'�����T���>?_:��\	�]�?=	<����㼑�>�>�γ>;x�����U"[>����� %<��>�p �|�>Cd=�g����:��>�*�=X����׾�d<��=�͹>~2�=\�
?W��>��J>��>�;�Z��>�%>�B��>���Б�V��=���>�"������>��>��&�(�;��~����h���1�l*���h&>*�g��!>��>?J?N`=>��=d�i=�m+?��(�u��=����׾�F?����	����I��h���A���0��T����>k���9&����>c�>�|��?i�g����E��链���<��]�~&��F��=�/> Y�>�뫽���>x%W>D��>��]ּ.Z,��fݼmez�s?���þ ��=�W����<� �>��=6N�>��������mm?�5�J��>���>w>�8V����>���鳂>�@ ���3>�?ͭf>M�C��%�>~ۃ=�,��$�9�?��A=Y���D>
!?��V=Ȩ�H���1S�>b�>��>Ҷ��E
?��>y�J����>� ��޷	�[�>r����O>Q6�>�����/>rW>p[D��N��u3�{�.��M���Ⱦ�\��S��>a�?BǾV�A?Bj�ߌm=�����d??��������?�q)>�Ε�,�#=��>�#d>|��>�Sb�t��?-�O?-	,>���{�>bE�nu����1
���nK�/��>���V�>�V�>A��=�z> �=��=�Ɛ>!�H�u����$8��T���H^��>]6^�:�`��쿾˵����>�L>��>����?^W�>xO>��\��Y���������=�t�Z-����>0y��� �=�n+>RB�>��=�}/�R�?��u>���>E�P��M�>�6���?�/W����<b�^>��>m��;�J���U�U��>�a?��K?6m��q�>7�����G���>6F ������q����⋐>=Q>y��<=?�_����A>-3��Zݾ>%�>W�~�U������>?E">�>/��͉>.� �l���G�p>+�?��?�I�K;H��:�ui?��=�;��_��>���>F$?�t?�ϔ�>|���v9?�G���ڱ>��=֋��05?��l�u��>��!?��B?Y��b?�i�>�$޾W[v>��>�|�=�!�=�K��%�<:�$>�^c?�1��Vt��,���ҟ���s<�24�R���x���=��7�%���>�+>$[o>�=˾�\�>��?��"?�;$���$��vL=|�>��J��;���Ľ�?S<�>R�_>e���I�=U��>�
)?J��?'rҾS�[�ev�<�`{>�Z;�3忾��b>hb>>��ھ�������n1>�xo�������7?R�={;d�!�G>D?�>
?_��>Y�=��ܾ��>&�׾-�;��.1���d?bg���H��D���>�`��B�|�V-%?�>,ƾ+��<�㗠>g��|� >�!?�<<z�>q��>�$�(�~=��M>܌%�L����L��2��n%�������	��>�|!�%n4�h)<mNb��iQ�r}�X6��*��ƕ=3c��������	?�X��$>�Xq?Ҩ;�n5����{�l?)X���5پ�-�9�>n���\,=z��>�<�>qо��n���z����8?�x-��������>.w�>K�ܽ.ݭ�=G�=�X<>��>3׾�?uf�<�V�_�>�-�>[,*>�s=0>O?d�ɾ{�e>�	��]V��W0=��= ��s4p���:��	վ� �e{�>:���ݤ>���>�o?�Z�T6�>��x?�׾��=�O�=B���U���w�;����@�2���6����=>�}��̑�~��@��>,�ܾ�=�>ŀG��	�>�"@�+��	?gH&�5D==r�4=]�y�f8�*��$�L>�w�yv>m=Q>����5����>Ŏ]>nN��'S�=
�>W�1>�!=�d�>��?�⼒�v?@)����B?�?�TH=�w�>K�̾%�۽�˯�.O�>H'I��v?��>�$���c?���>!?;%s>u�ʽ��>���Z�>s���0E�<)��=A��y�>Ǉ�<ڎ��ы=7��:X=s���P���#��>��|�n�p�d�[��!�=F���Ƚ� ʾ"��=a�$�ž��	���q6<�L����c?�i��]�>	V�=��D>y.�>I�/> �s=%R?	^3>�e?E�n=��/>7#?N�9�mK�>����gF�Fׄ>��<��J�/#G��?�?��;'�>�?����y�X3�>����P^?Lu|�S/�?�����>�.#���j�x��=�W���X�ԓ�l�>��U?������	8�R�
?�9�=��o?*�b?�?��?�gb?S�,ۛ�7��R瑽��=�?�s�#_"�-۾�:?dUJ���M?�,�l�>L$@?]�̾I�W?���>�H�?�ݾY�ÿ������- ������I&����!�?3��>,h>�VJ>G�q�>z4���aſ�Q>��>9�-�D�>d�L�f���?đ��?��g?Ш=���i`�?�>H�U�!��U?��R�T��ڜ=��G=�>��*>�����9�?i���A6?��׾B�Q�0"?���?�(�s:t?zA�?qK��?���+�>O�>��/�?��?�sN�=��n?̹�?@�=}�>r!J?^��>���> ���j4��W�hw��P�?5�(>P������a��Wt/?v)a�ֻ����^?ju������[�ᾎ͆?�䊾�*@�;��P��>���U�>�ӿ<����&�>.iϾ>�F����>�俥�e��ɜ�� >?�->�"��Z�2?�����^���|��@�?��I�rF?Ҋ��Z���0��>�ijF�#֒>K�>`i����V?$p�>� ��1���>���6K?�b�>�a��L
ѿrn�Ზ���S�T�u>��Ѿ�G�?>�������P
@��>��>�3�?�x3���=r�?`O,?�� >��@
b��쪿.���F��J��!�?0 ����=z��?��?������x�r*D=`.a>B���+,@7M�?�
&?��>	�W���?��)����Fd@���KD�_酾�]��`��d�E�JF�>X��?/�?�P�>�?�f�ÿȎ�?��̾����!dX?��/>�?�&����*��S.���
ھ������i>��|��\?i����?��-�&�.���?�,�>E����^=$(��7�����?M��^+�=��-?�¾���>��?� �'�"T࿿z�>p����!���T�>hc��Ю�?[T.>#�?�~?�-?l?��M[?�4����p>Dm���2�[:���\q>��I?o`�� �b�?KE�ص�ªF>&��>́��v���=�3�?��q�����@�=��*{��br?3Q	@�9�/�����?3Y>�(��Q��[]?!���͆��?�>ǉ?�t�?)�V?��-��<��w�?����=��w��m�⿆ӱ=���>L�;�	@S~�f �ur���Jd�2���h��2��?���?����G����?��B?8/鿒�8>#�龱q̾̏C�z����>��t>�Y�*���a\�?L�>?{�?F4e�!Yo?Vt�?�ŏ���=�Q<���ؾIi�<m{;��q���i�ʾ�^���#�E�����x��ێ��jĿ���?�u�>~?�D�>J�*?���?yo<�j�>���T�?B��?�?n_U�%����b�?F��4���1�G)?���>ݩ�>���=��>}3@���>F�/?*B-�ۇV?�G>?*o|�Aڌ?K�����?f�=!�?Q�{�̐P?cEɿA^E?�����߉�_�U?VF�?S|?a�o��	���n���4�;ȹ=�p��!�H?	�E�*�1>9�K����={+3@��7���3���N>M�->I����#�?�ɪ�iD˿�L\?]]?�-�t��E�?R#�����O�>��?�(�#�	@gD�Zh�>a�?)��?f#Ծ!���Ff?p�&>:�/��)��Ԝ?wvK?��D���)��?"�?���<iY��X����羭V>8z�ǌ>?�f>��?wh�?[?�Y�z���dS7>�����>�^�?ލ�?9������>�W@��F?s��;�ü�[�����gn��&��x!�Ү%?�� ���A?A�?�i�?�4��B��D�R?Ͻ?pz���1v�QX">ѻ�?C�e�	�?�E����a�?s8���=R��F�?�U�m[t�������?�?�`���(�Ok?�����)��a�x�پ�Ra?�����A?��Ŀ��n���(�i�u�5�'�E5���й?s?�ݗ����>H����_�>E��1?���>��2?�k��z����>o�?���i��>j�?aL;����*@��A�G��ɝ�>C�����о8��?����ym��=L@�p�?�#��ո<��=��cj��O���@��;�y����]>hWU>e������>b�w��zS?���>�XZ>=Rf�0=�?��_���?������������A>}��ｰ�l�>#��:����*��ρ����>[�k>lHa�����JJ��f��1��7H?�o����?�?=�d��с���@��$�#T��	�P���=<?i���X�>1Z?�jg?
�ڽ�Bξ�h@��>��S�5V��i8�=D>��L�'�����?���>�X_?�U?�Y[�5���?�s�?�;(@���<5�>Ȑ��ք?�����n���?�������1U�UAo�sH��h㡾��&�?&�߿)k�>�?��J?����z��2�@;|�)��?�Ͳ�BD𾂱?�ᐿK>��x�>*�����/��*Q��q�=�Q�s�?�S>�0�>+�G>a�>��n�Or��]�0�k�?��I������Q>�������s�>��t�v�?CJ�=ps����),(?�r��p����>n1�<T_������U�ϿP0@���=_��F��?�ʁ�`�ds�0���`(�>�8?�ys�Af�?<��?3m>��8>�L��-�>�y�>�����^>6̩�����O��]����2����?��?`f�?�c����= k7?MM?��^��<��Vb?��?,�?��)@�;{?�ۖ����<$"��FtM��h��c�4�=��h?xwÿ1
�>H��*�?�3ŽġE?N��?�돿�}o����&�`�_ ���=T���x��?�����I?�LI�
�4�c�3�8�Q?ˋo=~������]�?:.d=[�G��<��T�?����xj�8!]��v4�'����j?C�+��?眞>�.�?N��?�1��-0��M@��D��Е>AN�?Q��?�@'@�Y4�Fo�}`?U�.?�P�?�.L>��;��9�=�&C?T��?��{���ľ�ִ?1����a>jr�?�5��ԡ��!�?�N�? �����1?أ$��K�>B蘾b��>���נ�=\��� �؏��O, ���>�;���$�>�T��A����k>��>Fհ�6т�:�˿���>�,o>e�����?S����d>�B�4���{��>Q{/?�:Կc�Ŀ��)>cvW�e��>�����?<�g�i: ���>��>D4�?^}�
�g���;>%qf?�����>FT?d��?(�=[3�>���?��?���t�*���!?&���4*i�:(��#�U��?��>��=FI̽??�ݥ?�-�$��=����q�<,Й��:�>��SW�<�����3=���a����a����l?�(�='���b�#��z�>GD]�,���B����ƿ�����ˇ��6�=�!������1X?��>���`���^=~=���1�?�ޒ�@}��!lu��uy��e�?s�7������ſ[% @A/9?{�m��A��W>E�>-�E�۫�=H�?�1)��O��=D��;��>��?�턿8!�>��7?�o�+9E>l��/����s�n?���>B>y/>���O�B</�@�_�>�˫����=���>���?%z�?36[?L�X�j�)@�,?�z>m�-��X?B�>����-�?�2?��\�.��"�����ؽ���s�~>^ ���"�>�սK��>�3��5N�8>�q��^���-ȿ<�?��!�V���h���=o_���M����=��>�x��ï?�jy��Ꮏ����?�?::?����/A9?��ۿٌ�H�>K$����?B?�4�{����?�]D?%�/�ܿݳ?� 2���־�`�L@<?Q�!?�2�>E�D?1Z1�,���0c?��� ���X �>	i�����>QP��NG��9�L�����,�A��r>Uo�|,�
�(��$�=�~�>*�?���>~Rk=V�����{4L>U�پ��]?��]?ч��cv?%�=�IC<��7?�}��xc>���>sm�>��>�I�>V|>���=��!?]��=��}�->ɭӾ����OH�5���>����c?R��>���1c�/�=��о�=��4���x��=�e?ѡ���4���g�>~^���>ن=$�t>w��N�F���}]>�B��$,���}��uc��k�S�cǛ�uE�>G m�˓�>�����8?�4�>jG־M�$>�P�>��w>d��=`���!��Q�[=�'?3�=m�Y�g?%H��+��>1���y�4�L>���>Uk�<:YE>ۮ�>@�������qM`��ɫ�� ��L{$���USq?�Ǿ�
����L�Rs����>8+h��S��6v>=O�>�-q�:F����>?�>��>B�>���;�����������֋�;�i>�M�<q�d�k�/?��ξ�� ����uӛ>t1
�r�(D��#�(��~v>Gy����M�>�%�>H0�=C�!=SL�>%;��5���Nýc8�=֩�ʘ>����2A=��!�	�����1���w>ŕ���_�����Cy��v�$�}��ck�=��<�I>fj>�����y?�Q���=Ru�>�kżo��=��> �þʇ�>v�`>��6>H4ھ��޾��=tؾ���>*ջ�dG?��K>��R��Z�ɳ2��&+��-�>e���J�.���z>�?5o�>&~}���k?8��>��c�aF!?���>I���l%�;�R��m��2�?{�>�E����$>͆�;�xν������>e��>�"��W�-=C�n>�౾L�N�����˾��^>X6���;�z7�=Ps?��K?��>Y�>�Fj�������B?P�X��U?w��`��Y9���J��-��yz�69?<�>vl=��������>@'�=�B?
su�Px
?�M�=�8��F�2���-?ϯݾ"H?kܭ>��d���!�+��.߂>:��+�	�jF-����N];Zp�>����Ek�iaZ>V�"�>M��s�=$$��@�k�'��<>�/?�e����[��>��׽����?��8?P���3y��.O�>�ҋ>{7>�+��)��79�c�>Aʯ��N?�=�S> �>˷4�+!���o> �>�І������l�=˙>#"o>=?#b@�.�#?�.��,>��^�8~�'�=(v	?�3��j7�<l�9>A��>�j>�6<3!���k ������ܽE2��Wj?bl��3�Xm�=�K>9�?�d?��|����>-p)?��4�����(�y">�d�u�?�N��$��r3�=7Տ�AX��zi�<YЪ���*��[=�1�>�6P>�i?�y?D�>;��>5ž��<���G���7 >�'�;�D>;f�<fCj��e�>��?��`�?�`�>æ?�fq��v�>�ĺ>8����>��F>����~�>�!�?�1)���>PXe>l>�>$�����>�v �G,���͉���d�_�����㾂�>�뀾��$_">�����j?r%z?e���kN�>�p�<�_X?g�	���Q�e�>pH�>��S>!�	?�l���o⽶�߼�n�(��}ҽӯ��^&=>�Yž/1�><�x��v���<h�S��z">�Ʋ�H����o?<�J?:��h��>ϰ�>��>�ڊ����>SH����|����>��!Y�>98=�G�>���൯�a��j�f>�6���2��Ph��5�4?�Ε=�F>��,?�ž���>Nd�ئ	�-y?���=�R����U���>�<����=�K�<+���_���'�B�׾�z�O�b>�4�u��|=5}�'=b�)e�NbQ��W>*�)?8����9�P��=bz�>b�<��h]=�h��o��������Z0=+7k�_?�>�%ƼP�߾6tE����?XD�.w���w>�S8?���=/���u^���Ǽ��=�>K@=.Q�����1��}#?X�V=����4�=�D�>��H>�~�f�a�ݵ�>B��H'�(�L>ݛ�d#���tm�.�j�j�<���>~�>��8��x=�0?D=,�x�==��?��"��>(�=�G=KŨ�򘪽��?�z+���K���=w��NŽ�JϾ�Ž9?�>ˆ���m�=I1��U�>/��>�9>��>�:?�I�H�/�	��>&`�=e�<�I����3?Kh˾��
�����6�ݽ�X%=�b�Cp���>�����U���Yt> ,��/7��(�>H%��M�y��@}>m;=���>� �>�CI�q����+�>�*>Z������O$޽�a�>��>�_��g�>>��>��>��}�.?֕=� �=8��3)��/���Zݼ��&�.i#��=~��>��s�����8�>.!>�QP��?�r�>��>��n>v��>�?��W>��&��_���+?w;ۀ�D��6��&*�<�,1?�s>7[}���<?��>g,��}(T�p�ɽ�,;����ަ�Q���Ra���������3j�>c�=>�i��L�>'���V|���>�Gv?����Z�>��
?�)?��,�~l�>Rc�=$���!�>&H��F�	>3�m��^�>i =�u>�
��~��fP��ɾ��>)Ni����>�4����^R�>G��խ%?��>�����2��">g��c��ё��L�� ?#�?E��>��>�\�>��>%M��-�|>��N�}���Y�<b��+CE� >��>hX�>�-�>ɰ>[$>*G?Yf��f?��<�e?��ӾT�>�<@>d�>�e?T�?DM��c{�F���˽ս�S9?>����>�Ž�Z �d1�>������<���=���>���E�m���ѽ�2ھ��ﾒ�3�r�,���=/	�>�5w=��>�F��g�<6���I?������O�[=�6���+�N2'�Aΐ�F��S=�>Ƅ�
����>n�6>��>�*�>	
'<��L?"�=>��!�`�X��/U��_�=O��7_��KȾ���=�����v>woƾg���u�>��<?r���K�>�>�i�>�̽{3?�*�=-XE��i(�}�*>�?Ծ�d}�6�)?�X	?sߐ�ҹ>�I���g2?�Y�>����P��m��G�GԾ���>���v�> �r�җa>���=�����5���9�V�����*���!���J�}�����w>ižn���}w"�������>Ry����½J�>�$^�G`�>Ӷ(?�	�� ��M�6=<i"?n�����
�<A[-��r���w>��?��W����=�^<>��>�-?�����[����(<���-�S�۾�NH��>�Lg>�d��^b���>��C?������>n�$?�"�>�C�"1�=��ý�X�=f�>�<���>�u���>�%�=AϾ�R�鶘�T3�R)���N�P=�X�4�6�ݩt>h��3���>�V&�+���S#�>H���\V���$��D�G'A�����*P�e��s���J�=���>̒����%>�\?��`�IX��B��>B�=�;徙�>=7�=v}ݾ2�>��>;��oO>�A�>W�����h=[�h����>f5;���r���R=���	�|������>B�þ�b>�>0�>�6�>�_�>l��>���eI�>`�>>�����!?�Z��|7�;!��)>,��qݽ�.>D�5>�.�=m�S����<��7=跾`�A�\F�>�����^Ⱦ��<��5�� �h�5>�@�<�bm>z5ƾ�
�>�������-A�=��*��^�U_z>%>���2�ӏ��4��="��νܴ==�a�4y>���\����+�>��=��;��D��é����>�9?�qb���=,ӽ�v-?�)8��"�����>�LV>	�+<hʼ����>wu��ul>������0�=��>�X���~���H�4,_>��G>߯��~�u�)>��̾hȾH��f����E����P�����,w�z�������_W�	?�|T>U~�*?�|�>�mҽ��=*[?��>DVf>o�V�?�_?���>ޕ�=�����S<���>L����?彟=.�5=���>� �=q�B��>��m=f?�a�>����WC��a���%���=?���&���H��>�R���F<_�B���=�wھ�fW��?c���V��u>ʏ޾S7?M�9?
?3��=�B�	t#=w�%�����+��%�=�-�%�	=6"�\�>G�����ս�� >wP?��Q?�#�>�:���4?)l	>��=����z�>�ٌ����>|�1�
?��>�x��-�>��I?� Y>Iȕ> k@?�k�=�>=���>qZ��8���(��CL>0;>}q�&eؾ��9�.��������6��rI��S�;�c
�.�rO�=��6>)r������Ѿ)K�>��>��?�?Ͼʗ㽨������>�
��U�=Q������f�k����h�<����/>�|�=�l>
|\>E��
0�>bc?�c���V��^Q��Z->S���ߗ>A����(?��V>1&;��ȍI��5�Ō�j�@�!�X�ȧu��!?�-Z�Q���x���0�Jj8���H���ɾ��>�Ĺ�%<>F:���=eM�D���>g�=����"�>X�+�{ؤ=����d?�D����?�*��P�w�ri�P�f>d���;��l�f>�a�Rf>�$j�p�q>�����/�=٪�	��>_�?��>���>a��>���>^dk>=v�=��%?�y��6�>�ɾ�� ��Q;f����n>���^Ɣ>r��)>6`ӽ��>�����G��n!�{)�V@b=��2��x�?`'�<�n�<�	k���m>��>��Q>��>���?�ز�s5K�z��>�:��>��=�E�=hk�d��L���,B��mAֽ7�E?D�b?1���H9�>MC�<A���F6��n;ݼ�	'?L�>�J�>W��>�lI�>P�q�%>Bφ��>���=[ꕾ����9�����O���= �#c������C�=�+o=��X=0s=C]>n-�>C'�;�> �a?�����>{W� 5�?��O���?{����O<=�>)��p���m>d������1/ݽM0_���?�����-�=ǠC��d�?������>�<�j�>K�?Xgֽ*��?�(�?��t�[I�>�"x?F�{�}�>$�����>�#�_��>P8<�z�>Z�ʾ;�����\��j/!�������?�%�>�������t콚�[?s�)��<xx�=z�?u�5��V��,4=��a�~Ng�D��=�����W��Q>�鞾i#�=����OP?}�'>�q>�	��G>�D>�2?��E?�wz?�|��V��>䚽�@��v�}>��9\?�N?d��>uo�>Z;,�/?uz�=�!�>�Y�AF=��<?%T�>�S��j=��4=�U>��^>���=�� ��J�>�P�>�w�>s������ƽ<�P?�?<_"�w�C>���@I����@?v��(=?�
?[zu>��X2?
U�=᧱=�ܞ��A��@h#?Uo/>�Z�>3��lK�>��)��~�>퟾����=�u����1���>�4�8��>2G?m�>F��>Y?pΊ>���=�!?E�>-�A?�I��"�����W>��Y>g�	��_�����=�x�>�y�>�N�=P���m�
��!���I�Z]�hZO��\�=O �=:��ݩ0��q�>1�4>Q�t��\>���>+�㺹��-I?�hN�� ?�t>�W?|!���a���>.;?�G>��s���Ƚ��e��Yﾍ�5�:Bg��M�:sd�>�B=2e��?1�D�o�V>��=��!?#����q��#q>3[��C�\�m>Y�U������k?<J���ƭ��i0h>�$��M�<jE��g��=�D>� ��.�>"g>)A�PB��d��g�b�T{ývqe�_�>Ƿb=ߺ�����n�>�)��]#b���=�� ��Й�,A��Ap����>�#�'��]��;��>:��-#6>�#�xjM?��ż2������=�oH��)�黻�V��>���>�?�Ϟ<�|N>�L�>n�<����>
;<א�>�6O����W����6���#=�M>̥�沢>��>pk@?>�=�o�hϾ�{�>;���3>6e���?�>�����T>u�U=�x��C��l=gdL�3[�>�)�7�$u6�y�
�p�e>�|�4�����p�L
 ����>�?��_���<���??BN�Jbʽ~Y�(��>�'�>C�ڼb�Z�}�?g�a>k�,>��;��?Y\�>����C¾� �=b὾D/�7�D�M4�> �پ��Y���
�
��=a0&?�փ�R�+?*M�>�>%޺AkV<�������O&>�^׼��=�}n��O޾<�&���e?���,�����>���(�h>�Ž���?h�G�qr9?/�>a%A>&�>� Bּ#�>8&�>�R�>�*��#���:��(�*_�=Q>o?|>Wu�=���=߸�=wo�>l`>FH�����>���>Q��=υ��(�>�U>]�H>��= G7��BQ���%�Z�X>r=�=
�S���?�~�K�������"���ݾ~G8��[^>�b�?��=(/�~)�Vw�>)���v >��g�< q?��K�f���eN����?���>��5>�r�=/?*-�>�΍��� �v�Լ�5�>eӏ=��þ3�?��0>�=Cs�I�>G�Y?�#9?��?��?��>��r>���mY�?�5��O�B?��=N�A���)?3�>��?�n޾�0A>t�>������@��=��=����>f!=��Aa>yX��A�e=`(���,f=�f�OX?��V>��־�yC>.=��`�$>� ?�O�=���)A>>ń<� ������|#>�Ӈ����>Z���8�W>"������J���t?T�>`��ʖ>��:����>���>��۽��ý��k=V��=���>p2�>�F>^�*�q��>�哾 ^>�7?�ɱ>�~>`�>�]�>g�`?.衻��B�J3>�&Q>!R%����M�>�V>�o">�\ �X��>�΅><|�:y�=Kʾ�<�?����?w=T�� �o>jDݾcA"���?>�4&>�����Z�i�ܾ�g��Xg��A��P����<�XȽđ�D]�#�=�)%>;\���# ��坾V��1����	=vx&���*���/Ӫ=�fj��נ�%򈾽��>��I?
��v6>�0������P	�Y�>���>-~�2Q>06����?]�=��|=v�v�b>�>+�ʾ�*m��i�>���>aQ]�;YU��h��3�>��>���=�E(���*?���=�>��T??(>tu�<�y�h�=�yH��	���,������$о�q4�a����FZ�J�b�L�=�tv>�훾��G����='� ��	Ѿ������md��� �{+�	��=-�*���#��ܕ9=�[3��g��V��r�����=��ľU�>���{m�>�Ϋ���K�x{�>Gg��o�~�	*��1^?jo!����>o�_�]9> #?����&�w?-}?���hE��s��D����� �����]�ip�=�x>4��d���r����1+�>uw>�?�=?�<A�D��>�?�ޚ=ɠ>Y��J���2?:l>%�I>���>�j?Z�Ջ��.�;�{��=�x���>m,޽��>r6A�ꤾ'����>��7<.��=�s��?�S>���ӳ��v�^�?<���'f>��9�������ya�5���ӕ�����|#��ᄾ�{>>B��i�<�(ʾ]�.��򠾀"���/��sR>#��>��E��
���?$/-�T�j?�7b���=|�Ľ�����g���S������'��!?.��ܡ�H���ֽ��U��5�>��>���=N��>Ҳݾ4}[>8j�T¼e9D<h�<9%=s�=�U�YTo���Y�,�!�����,�����缞2����X���b<�!!;UW=�}=�=op�=b�=-�<�>��=N*=x{=���=��l=8̭<���<�|q=s�<��=L�x=E��`h%=�}�=�r�=>�=�σ=��>��#=�@=�b��4��TZ�~��I�,<T֑<�=N�=æ�=�.��;�d��8=*������p�<W��<��Ӽ�v1�Y�=�'�������=���=Gf̼�؛;g�=�zw<O����
x��=OԼ�\y��S��G])��	>A�=91>ȼ�=�L�=@�"=t�p�r�<�7�=jN�:��s���G6�=���<������;�=�6;�����&�:�<��=���=Q/=W3�[>W��=��=O��K����������;����o!�'8�g�I=�\ڼ_�������w�<�����I;��0⽽*=�=Uk�=J/={��=dy��Kj�ȃ��QS�<qK��d�:��N��I�(=��ɽV͉��7Խy*�Oi�=QH3=��S=ڼZ��7�:hٽ 䵽\����������#���ZO�I�6���=!st�����l<��]��U���Q�A�d��s��k��{�=�����g��&p�������r�������=�Ԓ���#��an�g���^w��V����K<&O^�eo�=e�=)�¹�����>�3�=��<7|��>��*�;�-?����=�=F�.=1A�=���=HZ��𞽐L���z=t�$�0��wź�=�A�;��@�Ǡ,=��S��٪=��<7�=�=�s���-h�vz6=F���#WU��{��U��=���=��;N�<������=5��:�G�=���=%g�=�dh����<a�n]=�=�t ��T��<��=�T==�厽n��=��=��=%Qe=�M�<}ݻ�}=�}=�.T=e�F��U;O���Z��>��vܽ�-�,D���?T����;1[;�D.=���`=�ľ=���=�<�ض=D&>���=����ƾ;^�<��:?�ռ��~��ٛ<�������5����2���.;�F���3;O陼:eH�����լ�=���=�=h=jA�)/�:����=�܀=$��=��^�%��<�d�=:"�=Y�M�ݧ�=��=(c/=H�Ž~;��Z�?�=]�=;�L����' �/B�=��9Gl��/���=0�<�v2=I�d<j�>��'=F�����;�^O��}���.�<i�$<��<S���F�Q=]K�<�l���%(<�	��'�v<�[X�hl���;c�����zH�<\]�=� �=�������=��=��=���{�����;&�j�9�۽)�=>�<2v<=�n�=�E����>�xwҽ���<~m�<�+˽�C����<C&�=`=\qg���=3���fͽ������*��pD�:�=�=o=�|�=��=��=��(�`���>!�<�6�<�=.�`����<�+=�X�<�Ӽ��!=�(�=[aP=ւݼTC)>�k,>�ٵ=��Ǽ�9>i9>3�z=�C���	q��y<(+<��;��R;� �:���=�=�uU=Ƽ>�J(=B�v<�Y+�n4�<�ٳ��-�=�%�=B�t=��=���6(�=��=�9�=Sw=L�C�d�!��(@���M�P���e��<6�=�_߽�rc���8=ѼSՈ��H�=&K�=�==����=C��=��
=I�Ƽ#�>�W>�
\=y�=��6��H��^�=���=c&�����pԼ�Ȥ=ۿϽ̨���>��ː�;H��E������<�Ȭ���ʻ=��m�ͽ�=��=�Ny=B%U�2��=�k3>�y=��Ͻ���%Q��H�i����	����N��̓�ɔ��ǔW=A��c\t��}�<H��=������w��?;=�m=9�==�f��a��4U��ߨ���"�4q�z�X�T@��܃<򟌽��w�ɪ��[E=�,*=|b�<�qz��qI<��=�E��=����B�t
�<Rb=ItG�8���^�9�`�=W���^����;H����Y=�ۼ�0�ս2�d�t*�ъ���,=Po���н�2�<p�>Yt�ԲF��� ��(�<��:<���$d�=Ӏ�=1N����	�R���֛���<������=�%�=h-�=t�}��|��g��hK�f�̽�d�=�#=����̻4�=܁G��ȻEL��_[�=��%��!����޽�>�=���� ����׽�%�;��:Z���9t���s����=�]�<��o�T�)��9:P�<�I�ZG���i����b�=��
<>	�=X�=Gi�<���� �����=���=m��;��{�V=�b<�(�
���;��=�}B<>)���E̻q�'=2��=�[!=7J���"�� Z��J��q溽�p��k#>=�I׼7O�,��=��Q�m��=��=�W=�[�w��̦=r��=j���%�b=��<��=�h��B��P�{������ˆ=��F<��=��D���,��=|^�=���<h��=o�;��l������߽��%������9��A��<˒�=�:S=�U��_Q=�>�;=Fx��d��=�c��#�=w��7�=59�=�L=Y�<�ʪ���I����f�<f`�����/���'l��A�����u_�`6�RO��JK�=}��=���<>�.=���=�DJ;]�F������
=�Q�=�i��k۽��<�#�=Ť��*ǽ�}v=Gp�<;�ս����H�2�!���ȼH���޻������C^�QK�=x~>EE>��>e�=��G=صu<_��=W��=uS�<�YT��-+=:�=Tl<��&3=\�N=���<B�<B�9l^�T�C=��+<�?~���ý�}R;EQP=1s�=ꛜ�	(E=�=q=S*�=>����5��{Y���n��;���H�1��=B
�=�`���=�&=ٺ�=+7n�z�?<�B�<wL�=�����p�ؐ�=5�=h��<���=�̃<��X<�)�<�4�<�.�=�=�3n�N��=���=	@�y��ζ��m�W;;�����ƽ<�^���*<�������=�>L��<��#��x�=��=Kb�=�7=>�'>*��=O�b=��׽1t\����LOA�+۝��+i<沍=V���i�$��=��=�<t�~�]��=�;>��s�T �<�5n=�3=�� =(G=��������<d��w䃽�&=���Y�a�� '�8�+�Т��-���a&��0ν�{ٽ��R=����Ce:������F`=eF@��1<6�����`�r#�=� ���½[*���ꆽ�락�|�X��<���=��n̽�1�=�G=�1�y�v<L��=p�=�(����;�.Q=�5=�wf=�ɽQɡ=/��=�d�=���<�<#=�1=�/�=}�۽����U���1=�9{=��j<��¼)�7^�u=N|��������-:��:E����a)½4x��:�9����x�==n��2U<��=�{I������:����<��ѽ֐��5��d���*���꽇y�e4�� �~D7<��=��><0��!���=r�l;��A�uFԽa>�aK�޾}��C����=]Y�=a�:�4��`Y��T��<��}��8��L�=D���L�Yν��z;\�8�ύƽv�;;��=�[�=��=���=�7�=q���r�;��<��R=Ⱦ�;��ü���=��=�q�<�u������b�>h�;&�=�E;��=�e�x��-�����U=@0�<�+�G/��4��<JSj�7l�x�ܽ1��l7ӻ�[��+޼+Ο=F8�@�m��8��Duƽ
���X��������=�Ӣ�z�Խ�3ٽ+l<�cg���A�\��<<���j���_C�A�<�j=��½����E�=g(����<[H#=��ZŻ/h��L�9<�����<��;� �=�nF�F�ڍ�<V��=LVX��N��lO<���<�Ϳ>yx!�������Uw�=��=S�7��sA�>�S����W���J��P�>��o�2��o�l����0�8����⾈W?��?R�G>�Ȗ?T�����\?�>�1=��>O-�>�����R���E�Y����=����f=�>���>�3>$�>���=���>j�	>jk��a	��[����ؾ�Xi>z��>�qq��N2>�s(�X���&�!�F��M=��t��,��f;���>'%m����aҾ�C��n�V���� ��=,� ���=|2?�>N�<��*��+b>���>��7�{|�:oȽwQ.;F�]>�?{M}>���>�M߾�����Z�8��% �1�=���>y�
?s�>*��b��=�������!t��� �X�d��z�=���>h,?���=���>�Ñ>��=�u^������ߏ��i����Ϛ1>5L꽫㫾W�l���Q?�~>jܞ�Z����}=�B��I:�=PX�pr�>�j�=>��=r����%,?@!�>6��=\>}N*>�TѾ���Qj����>�8+���t��j`��%�>�F=�K�=���׎�-�����`�������$><�>\?���>�1�>`������Ϥ��/慨�"�>��>�>���l����2>�Q�>)l���<c�V=޺��&M�3�x����>��<�����E)����ƽ�_��l�>�>A�>�3?e��>M���+�?�1 >oB�9�� �����u��x�
��ȭĽޙ{�!N�>
˔���@>�wO��<��32*>�RI=��
>��f��ұ>����<=�;��vO�>#F8?���>.��>��"�w�H���	���&����p� <�$n=|��>�8�>-�վE�n��b�=�,�_^	�6gT=�|�?j�������;�F��;����9�˝��s�<���>��<�?'�>��0���>!&4��;D=� ?���>�if�تf����m�R��ľI��=��F�Lְ>�!=���������z!^>ҼI�N=�o><��S?�ߣ>3L�?�=w�N?�l�>�R��@>)�[���!?*���N^���ҾiCܾ
�=U+C=q�/?�_�>��J��3���I�����Q��{�$!�3ʏ>��:?��n=XET>�S����>%�g���<�=~�><#><�:�*����>۽>2���`��X�$���s>�h>��>�ƾy��=w;ʽ��Ѿ+� �����-����=�1�:uY<b"U>�۽��><%�w�L�p(\�L�T�FU=���dԱ�QCj=�媽Nȼ#�ҾZ��<+�]>aa��K�neR��Z��)<�9�M�7>�/k�ϣ?�&�>�~�=�E�>;r>7J(>Rs��Ù�=���A�=(�^��b�U\>��D?�`X>�Ο�������<6���L���)[�&7^<_P>�Q��6�?�?[ȓ���
�ss ��;�<�>��?�a>�b>�l���W>zk���V���=w�?Ux�>HC�=Wj��5l>�ُ>�S�>A���m��/&?�߻T�н�Ӆ>���>P�M>���s��D�>�~?�ז�)��U{�/�[��S?9]�>g��>��M?�;���L�>�nK>�"M��!����>����=��6���=>Q��=��Y�ᬃ>H�.�,��;�H>�==)8��N��*��=�\��$�/N����@��K��>�=?t��>�d�(<��>�V@�q�g��Rr=���>�.=�����E>��>#Ll>��=���H9Ǿ�q���v�=J��=���1�>�^s=n����"��#��{��>Hxu�M�⼧��<X��>Y~��  �ى��8]?0�V>�D�>��>5�`?�w�>�E2���u��L=`�`�#�ھ0:��C ݽO�z�*���y��ܺ>�w�>i��>
Y(=�W�=�Oͽ��ս�{ݾ-��^#>S;ͼnWS>@��=q�6?f�m�"�e>Ϩ��=D�J���h�>�}�'���>�5�>�	����3�J�S>�?M�񆱾K�t�����h?U@�>�q�>�n˾�ib>3v��?Y��:3@�+�=ǹg>�w�=`S̾�����n^��Ak�&�aֳ>l�>�G�>Ļ�>M�>��B>�*$���ݾ��ʾ1�<��>*y?�,?���>�c?�5#?>��e�C�z���9��H���b���3����>a5�>`�&�|1>�� >?���>�蒽0�==\�j�F>AQ�rK����8?0�}= \��=����P?HG���"�>�������܏���ýQ۔�]/>�v?V
�>�
�F��'�&F(�u�f��dd�+�۽��ܺ�F��>6��>ǽO>2�?��Q��4����%�Y%?ONK9���>�M�>BQE>�]]> ����,=F�>�Z>O�>�<��Ǩ�=r|��m>o���ѽrD�=`����Ͻ�k�����>C<)���N�Rʒ��:�w��>��.=�9��э��L<C��= �����J�Y��(�>�)���žy���wľޣǾi~>��I��S��'X���"?E>�Y��ǮS>��??���=�l=�q�����G]i�׹e�Ws�,���B2/<Dsm?���>T���~���MJ?==#�)��u>t�?��>�0*� �g=�f�>l�?�vD�1��>�{��TcY>�}B<�'?똢>�y#��y><A=���۾N1�QE���~�>ɶ	>�Fh� ��=_8>jA>�m?��{w �g��3���+��<aT�=W����WW>W �>+⼕a�>��W>�9���->�}s��?K秽��G>����R`.��Dz�ӑľfM���&>�>�� ?x�>@�=���?=�=�?ލ�>f�����I��3����>7P�)8�>u�>�/?C�?���=Dbٽ�>�>����(�����`��?!�9�=j��>�DF=g[��Fz.?�u�=x
�s#׾0���D�9�9�Y�Qw.��b���2C�g�#>��U>+鲾[�$>z�(?�
+>��@�⽮�?��>7��1��乪�>�Y2�������>,�'5%?j��>��7?
;7��X?�=6��n��$���ھ��R������K�W����>��@?V��>��S���>u�X�����c���>�3>�z���>x�>G�m>|�.>ݭ�>���>i�i�s��gF��-ʽg|;��c#B�>�`��4�/��=.a��y�H�=�0�� ��E�=S�2>s����=-��>�$;��=���]����>�y��`Ͼ���c��z@@�9�������>�lZ>��>T�?��<=�¼��� �־�� �oQU��]���&>�C�>4��>�w>�xs��L�>br���i�xn�=�k���⇾����1�
>�n�>��0=�������&ܾ-y�=Ƈ>������E6>�AB?Q�\?��SR2>gO�?"}�>sV�3�M=ڈ�W�ؼ(>�5�U<T����}'>��L>]��ͧ{>|�>��컬�����.��`?��w�$D��C�s�SN�>2��=o8�MlS�=�Q>����)=%��>�+�d�طH���>B5.���0r����S=>(��>��(?�ɤ���4��Gg�vX.�aVQ���'�=��H?߯��"X�>�� �G���=e�>��R>ハ�#=ޚJ>��,��ꇿ�K�M~=Ϙ>�DE�vO�� ?dw����%>��=�p5?��Ӽ�I>D���e!,=��o������>NC?��>�E>�١>�?�%���˰��bz>���>p�پ� �35)�F�>Ǎ>��ξ�D>��?��>�2�=�˯���*?��~�U;�������e�Vm��OǾ���>f��>��7�~�\G`?*����Դ��ӣ�,��>�S��:پg�%���J�ߌq����q�E?�K;>���>n?�pr�Ph�=��W��N��<N��X0�>�#�<���B��>F�->)",�ҴS<���׷�'���65��{5��`W>!�]>�Z�>|�#�V��aQ�F�0>!h�>�f5=�#>P����5>������˽�\���=,̽��߾qa>/K4?���jy$>	����+=F��16�x��>~��GY��^��>�w>��?�J�>ԃ>�.� ?��>k37>
��G�b?�?>]6>Ս=-B,�*��ˈ>	?'�8�=�9�Y>�@�=h+޼]ʄ��w���>��x�hH�>O�	��(Y>jjx>o�>����8H��y^=>�f���q(��(�>,��>$�羆Ǒ>n;$��v}>P�x��"��&��>ݭ˽�H�놚<;=�> />g���P��rQ?V�Z��k�=�>F���?37�>��;��/>��?��q>��<(~f�l2�>ՠq<=�"�j���L?n>o�ܾ��{>�@�>A���
��>���D־ ��,�6>���>Nx =�	C�N{I>���>N��;
"����I��G�=�V>�o"�GAӽ��C���n�>�M�����<=jU��>�y������Z��le?ǽ�?�� ��YI>$,=D�>վr�>��������B��U�>��u���m�r�з+?�Ȩ>���>�ᐾ��j�->�'?�%_���ݾ��c=|��iR��/U�	�s>�Ȧ<��Ⱦ����½��+>�K�@[2>�d�=m�p���$����>��c�}��N��ey8��ћ�yK��=���P?<q�>mV�=���z���I�����ž�p��ؙ���b�>�(�>;x��i �9�M�E~�>&dK�wO'�ڸ'�������׼�>m�-�d�>��w= �N>�c�r�F��}�=}�>nԚ�4M(�� ?�ɨ>p/���>�*>��>+>�-�>���>s�=��.�^㿾�� �����z�d�y򽾊f�>K�>ʮ�)9> �,���f>BЉ�IQ4>��>��>�ʽ�vϾ��\>)4==X_�����L>�q�>x1?
S�>�~?]���z�	>�uվ�%G���j>`�d>>�cG�>?�]>�m �X��3ľ�(�Nʛ>���\��(߾�#��M�+e�>G���v�=y�?�d>\����>�UŻ i�>���X��;پa?Q+>��G��� ������9��2���yzڽYm�>䟌�����4��>M��s��?�>ղ��T��=ߤ�<y��>���>����wb�n��>�t�>O*�H��<?�_>�?����u�;n�\"�O����fW;1��j�a���%?�{���n�6 ؽZ��>��پs�,��2��>�RH?�mE>�6�>�j�>?�u����>��>�U|��#����>j�{=e���@�z5�=(>l�������<�>G>V��BǶ��Z��:������.2>-�j>o"��/Y��Ӄ>�MA>T୾�DҾ)
7����hU��;f>f�U����=ݦ>-�u>$�e��A�e1�>�/@>	_F����M١>���>�%?�s�>5�
?߰����F>��Ij�T����z=f*?��K>�yH>؊�>�Ts>|"Ƽ0�P�!=P����=�ҝ��9���n����>B�Ѿ���>5Oh>�@~>�[&���$>1��>�6>s��d���Q�Ւ?6W�8I�n�1��>��f�:�>G;�=6\y>��>�7�=�Li��k�A�?���uad?3Ä>���=6Q/�2$<���G�ؕ�>��M�q>&?*�>�����R���hK�B̕�H�a>�)��9�>�
��_:=���5��>�,g��>>�>ɏ�7C�9�>���>?�m�6پ��=壆�C��=�e�>�5(�O�7�
�O�D��>3��U�)��4#�Ç�>�]d���ྡྷ�a>L�>F_�=�' ={�-=�j�C"�>A&���q��dH��ս���>�p�����;��O>V�%?�j��2�2��<��
>�!�Z�Ҿ��>m�>��7ݾK�1����<V�L>X���l������>�>D�P�]�3�?ޞ������/W=���O��>;�7?}��������S���==p�����zо�8\<'A��?c�>Q�ƾ�B�>������1�z�]�T&ܾ|�����>6�>a����
<�k=ङ>��/�Pn���m�>�ٗ�o�bn�Pѱ=7b��f6����k�>e=!��ko��J=r�(>!�!>(�7�n�Q��?%�O���f������w>��<�O�<is�>�^=ޘ<�M��=���<�=��<�
>�[>M^A���=�6���&�>p��=�#?������(>́��Gξ�z��1c>(?��C�H���^R?k:����>� �g!��4��u�	���\��Z��0c�=�}׽��=�[6>�|��x>�=e���ݾ��˽��2���8�m?o3�֢�>�9"?�_S<L�F��Ѿ��>3��>�0���7�p�>�'��[[����&>)��?���>�O����b#���U>rwd���<�3FT=�[>JE]��I��9�>�d+>M"?�f�>WY�xT�>j'�>�i�A'>f��y�=:�	����������;�#c >۸E��[����O��-���J��@�_@?̤����!��%����0���>����]e�>��o>Z�?(��� �|T��z����rp=)-��'~%� ݝ���G?��u��d_>j��>a8�>3��*�>�A>ho�>�:�,�ؽ�i�Co!?�!>�ڗ��Z��}���������>UA<^��>q�>9�(����=�)��I{�����>2߾�>��u�>�Cc�r]>@��>��<�A��ܾiF�>�j1>R�����>�?�= 1�<�Ɖ�u[/?��>�⽱�"���,> �?$��}��;��=F��gҽj�1��o�>0{�=ɟ�= Z�>�j�����=]�>�>�>�U>7z>P�	�>¸����6?��;�[�3?d[1?��ĺ�>R�쾥�=���=��w=!v�"U�=�u�>�P�������:>f����]>/����{��`r�N��>�K�����>�B�_"���}�>}s��X�==Y7>R��>�n)�̡U>a߽pF%?��p�Y���:�Pwt?'üB��>C�<D���$g��[>\"?�گ�Qz��
�>E[�>1&\>�X�&M���e�>��a��}۾^ʘ�E\����]>�K��-�>+��>Ek��r�Ǿ�OE>Mi�>�eٻþ���=�x����>@H�)��<*yֽ;�A� �d�;E.>{��=&�̾|�C�v�r>R��>LMP�rx��x���e5R�����?p��=�k><ِ��p>`s¾CTѾ ~�=�G�>�I2��u�� �=��>u8i���W=�;��T�»;Cu��أ޾���a��<�ӽ�|��B�;����> ��>3�,���{9�>�N?��e�=�����>>�T�oGE��G��ؾ>�?F>�6���Ǳ�ӘO>vI?XM���w��g�>h�=����P���5@����=TY!?��㾓ʚ=S6?^+>,��SE?� >/u>j�����ȶR�D�O>���>"~�����=�ލ��m">J&���5��DM9�K�>��@��� �i4=$��>�+��J�=О��P?J��=COu>򝖾���>SU�����k4a��4>���@�$���=� �>�|���2+=�x����ٽ"к��e�6�I??�>o׀��d>W�>����=�<h�Ͼ'�>4܈=�'���N�x?�>�j߽������ɾ�>C&�j)�nW���>*>������=���>nVk>&T7=v��=A}�>=��>�:	?{��>�m�>T���-����XB=I>��>9X�>�>�?=k�PX�>`�>��>�!?a8?-E����=�����q<��?�ѽ�>�7ӻ1����E_��g�>������>1{;���>�l�=
 �=9�9�K�>>�;������󫀽@��>"6��:6[�������>+Z�=d�>�_5�CP��C�l?߽[~�7<ܽ%��>��>�^��ot�>-�i��͑�>4����>��>�C�)�q�)ȋ�d���-� ?�-C=�Α�v�)���N=��ϙE=��?��?ᨧ��������\��>f�>�h�a�=���> k#?ߕ����!�jb~�6��EY�z�߾�:ϾD�>���t2�&�g ����>��D���>��?]#f�N���WC�>N ?�Z ?f��>N�	?d^>��>#�>�Z=�,{?��?�7?�^�>i�5�6NԽ��=��>!g�>o��>��>�4J�*���pw���ȾWW&��OJ>�%�>���X?ý�>���=i%ڽl?�<��G8�x�I�F�l�>�"6�d ���k>{k�l�P>���>�~>k5��3%ƽ�b?���>H�������>�i�>�u����J��1�/zF>W#�>�@F?.�)>E*,?���>P�c>�d�=(2?���֡Ƚ_�W=Wc�=�T�=zFs�݆�K?Sg=��?;(0?C<F�dګ�n��=��>�T�K+v>��?;�
?'Ӕ�n�z������Pо������E�|��
_�=(O�>_�<�=	�J���|>}�Ͼa�C�(��[(?�	?±r=�%��L?�$ھSQh���ӽ���>���>��s��<��@?*#�=�`�g���5i�?,�*�B�/���)��&�c�^=<��9+���Ͼ'H>�3�Ln>@�ؽĚ��﮽� &�O�ג�u"/��*�cxO�5l!��礽rzC?�!<�X���ƥ<Ty�m�˾8C>�-H�	��?v6���`���6>0؆=N��>�/>Qy�=��w��a>h��t��>X+�<t@>�ҽ�0-�߃��ƾ�5���<I���KP ����>u�=1�Ҽ$@A�Q��>��پH��=��������:���:�=儠�)v>��?��d?���=f�?BHb�5�0�|Ỽ/��>3��E��_z������cK<�tؾJ�C>���j�������>sϪ�"sӼ��'�>?x���K���� f�>Qf>u�>[DS>S��>g�_�5q`��̗>3+�>�&?��>�`ھ�iI<���C������i����>��оfh�'�8��mؾJt�>m]\>����l�ݖ�=W�>�=>�����>*k>�<>.��+��<��?�q�?@)���5���B��8]�����?[<@��>�۩���վˑ=K�x��ϵ>��1��T��@�=�-��k?#0=�u��X���I�>������1>�g�L�>�W�>1T��\����1?aq6��8�>J=��nE��
����=R��>?jT=��z>���D{	?2�OR�5}>[�C>����CyE>�.!��ʢ>K[>�<%>o!�<���:=��}=��B>�T���D>%��>Ecg>��q}>_����k=N�\���>-�D>2�>�t{��Dֽ�f����>z6��cH?�j=�E�{������w��՞%=����y]G��E���!�>�����P>���o�>�S��6����0h�>^�>X+?��5>���>F������l�������>��>}�k���d��G?+�?��>
+?�#F>�v?�@(?5>V�̽�:�>GӬ>&L]<ͼq���?,��>E�$>B�>�{t>a1���>A$���+�>�x�>�sb=<F��;��?��������&�k�>^3�=��=�K�?���?Ce�>T6?t=$�k�>F?���d?�q�>���>�>x�=�>��?��v>\�K��H�Kz�=��=�Ծ[ѾU��=�}B��l�j�>]]�>�ܟ�c���K�S?=�K?�Z>�M׽y�h����>h�>�g���E?�+X?[�=�F��P���󒜾�0x>��=��peU��>�	���[e���z��2������Ũ��`d_=*�>��>wk�>Ya���䊾咽������꾣��?��>���=/;q��7-u�Í�4�?�������U�ǆ�����}�=3=XU�<&��z�'?͜�>U[�>qwM���>��>pb�>g�辑��>l��ƺ˾�	?m"�����=��P=2#�>>X��"-~�Vx��d�>{ک�I]s�����?��2��%оmR�������:�����=���	�P�>t��>��=�M�r!>�>:�=��.�������	�-X%�2XR��h���J�J&��� F?�G>�wŽ���F3���~H<���>ϳѾ��j?���>xx���v���%�*��>�/t�l;�'��>�ۊ����^у�%"��gi���]��>
?؝�;�Q'��N��LaN?����m~����U#'?�Z���q��P��=?�;=>��ؾ��w>���߂[�x�ڻ��Y��1�RF�=��
�e����O��	�ꒅ>3n���þ�羞�;���{~�>��>��T�Pt$?�h����
��QU�@9�>�S��i����1?��!�><Bͽ%n0>���<,�>�a=g� >��Mku>���>S��=Ͻ�ئ{>�-A��-�=:�ڄP���k������d>��>�O?���>^\�>9,���>6_(?<v�>�`���2>��>�'T=�׾t��.�nT�wF7?
�> .?�:�=Aa>؛�>J�5>�dc���?K4�>A*y<�r����9��5���d��?��eﾂl�>�/?-[�)4��{2?U?�4>�T��Bݽ��>t�x>ϛ����?�@?,�>����ƾ��>��|�X�<��>�q;>.��>��B������W�<�C�=���EF���,��)���=��N==?¾���>G'�<8�=+�оl's>�q��]�Z�Ǿ��(>eyx��w>�;>�e�>���l���˾=VW=�x?Q"�<[�ʾb�I<b1Ҽ�ާ�s��H�<� ?��\?}./><��>�o?��>s>)�=��=c��=m7>6�'���>�e���ؽ���4�>�����Y�>�I	?���>v �=�;�=E�:�[�ZYc>I^6?����P
�>͵�=R���Y��;�Ѿ��߾�gܾ�[�������|�>��?ܐ>씇����;(�>�՗>�p�����vI ?��>`Gȿ���� �bY�>�ð><�?��.?�M׻�|8>rO�>SW�>�N=����.J�>]�??ۦ=QY�ȼ��0�%���h=r����Ә>���>P��J6�1�3?ʁG?�M>������g$?���>h�;���>��N?د~>=����2>'�>�����<*�=�?�lǾ���<yB�>��V>�὘sO>�w�\h�=��ko.>\�'�[��q
>�j>���+7���_�7���=<%=���������>ғ¾b�f��ϽKx龪8&��R<g�?� ���侟 ��.��!��>���>�ʦ=��v>G9�w�=1�K>d̀�*3V���<��ڽIr����>v�>�GC?v�����>��>}��>����(?�)>���>��ڭ�R+?��=?�r�=jC���H1�sn�=�#4��S?~}?{+M>���-� �nhQ>O8>r~�>)��������=UӇ�A�,���h�
>�Ϣ�<Lq�=�h���Ҿrc>�= ��GS��V@���f>�L8�w�־���=�4?&b>������儾��ѽ���
��?�)�W�-��	�Z�6��ED��>�v�>�>d[	�$fڽi�>!�T��{�� b�>�5��P>�~=��8����>�ū=~�w�x��	�� >�S3�W����3"���U>N(*�CP���I����>���>Z�=��n>6Z?�?��>��?x�>�$>S@>[\�>���=�ַ���;<X��^��>񕾾��޾]�>5;�?��>�K>'>-�f>����I�E�_�Kާ?;�=�3��Ѐ��J��>�Z��������h'`�m׾����
�=oY%?���� ��.=�������;q�н�s�r�	?�����F��q;�u��pS�(/ʽb9����[��׻�{7���-�?���>O()=�XT<��>+�=)�v>yQ���'+?>C?y��>�<x�`�{��^)�uM�s�ži�W� UʾS�>��}�پP����[Ҿ7~*��Ϗ�v$?/й�D�S>(?�|.�(ׄ�xg���>��+�|�������P
����=��Ǿ��D�T�?��W?�?��D�����?vj?�?C5F?ɪ�?9�?x�,>>��>��[?k�?L>�>ň�>�k��*B?^L&�hˏ:�<?��=7!Q?�?�5?$<?Q��?W��>ǖ�m�>~g��v�Ӿn�M? �O?�e���\?�|�>e�/�#���k>���e��j��1��ǟ�w�f�ލ�=!r'>����ă�����E�>Ɍ���>?�h� �>?�0��Kݾ�f�E��>�{=�#�s"?+�?��:?=t�?َ�>Y�>x���.�>��C�ʭi>�D?�>�!!>s��>e`�>�?��?�%��>b�c�:���î?P��r�]>�4*?��?P�C��(v�O
?���>����&��a��ܤ��Ǽ������޿��N��>�=�MH?��	��ρ>� �������[����J��C�?��?�0�=[����P�=�==�{?熠>��?�`�y�Y�Ѿ7a�>��� '!>�I(�z�$��u���/>q�h3�.�b��Qھ_��	�@���>�S����<�����|ֽM����Ý�M�̾⋿6W^�kT=�͐<���aܾD������>���M(����������i]ҾD���ո?D�b?���>e�=��I�Q����9��m���.������>�q6>�2����t�>;Q��b���!�ؐ���Kc��ri>��<m��>���|(#?��?4U�4�¿A�C?���u߾\e/���=���Q?�>:ͧ<���=La~?��S?����i��>�$���þ��c����P�Ⱦ?�����>0��������
<N��־u��֩&�i���z�?6��>%��r��?"f)>�ʲ��'���N?���>$��<aq5?���>7����]?_�A?�@Q!��o`?$�>�Ӕ����?�����vU=�Ls�(�==g)W?�C?�𼝵�sX?�6?؍�[����{?,?A�?rj��?���<	�>��Ѿ�<G���=�T~�h�u�T�M��"Z�w�!�)�o��>?�쬼0�>q_��|�1;��K>�_�Ş�����>ȔG>��?0��>	0h?#!��N�>bBE�x��?��X��u-�t��>�w?��8�4zR>�~@>���U�]�2o7>�f�=��>9�M?�\��u�>��;��X?��?h}#��P����m?V=��h1?��?A�%>C:�=���;��c?e?�D�>1~��4�?[�O�q?�?�?\?N.����G>x�I?+�˾�&m>�~=��x�#��>=�B�v�J���cg?�jC�����*M0?d>�>\Cn���>�L�L}��Bt|>;ھ�Q�A�L��iI?"�?������Ô?��+��EA��b�y�>.}!?mE%?�@�?�>?`�=,O��	d?s�ȿ'&#?op3?�/�>�>.j�>�7i������6?� ?�>��>WS���[�?W� ?x�a?�O>Oe!�~�.?]@?�5���I��{!?�>L;�>�Y�\���>~�=�GR��?f�`�ZJ��M�>r}̼M�?���? r�>�f;����_�G?M'�<dMy�"T½��б�'BJ>D<�?[�ž����O?��?��?�'=-��T�������&)?�Ҋ?*m@?�w?�>g�E?��?D<*=E�� ��?��;?�j�����?-g�=��>pu@��9+>a�H?g,O?C9������	օ��ý=�-?�Oy�E'Ϳ�k?��=�t��n���=t��=�m$���꾽%����g���t��>��q���O?~X>���>�]>/�u>�d�>�>����6>*>��0��TQ� C�ݎ���@�=�괾_��>�)��5{?K����c5>C"�>ݭ� ��>LK�>5s�>�丯?6�X?�����{=�v
�Y��-�ҿ����w����������{������M��-����d?�cY�<ƾ�s ��d
?˛>w�>���?l����=�ϴ��,�>
c��*O?�:X?� ?����y�3���"�޾��P��OQ�%����N�?ca� �K�wĵ���S��}���V0��L��!>Xp���^v?l�B���>͞;?jR���{Ʌ��t�;���칄?�3�������i���Q��E�`p�>���?5����=�>��}?��e��m��Y�#���>�N�>t�>�7�X�
>�* >���qg���l��$���)=�׵��{��?��p�Bl��C����>�+�=����[��dH�Zׇ>��$��*>V?�DY���v>>�J��#ؾ��B�?�Y>�*x�p&��H��>.r ?u���g�q<�5�>U�w>#�h>�,ÿ�G2?w��>vS����i?���=�𞿝�!�9%<;��8�{;�>���>�FI=��i��֩?���>v�/�B���Ԓ�>�hm�ǃf?B��5�=}GK>h��> /b>`\���뎾�d���S	�B�?�Ͳ���F�eJ�>@3�>.!> ��>�%B>�Ͻx���̻ M�;�䐾����j?��+�?�̻?T?�Ⱥ���8?��>��> ���>��C��?Q3�=i�>=�߾>�GB?��:���ľ��?�y?�U7�f^�>R����8�>�-�>�Y߾�=I���=���<ꦊ>��i?��=?�֊>ȈM=�������?}|�>��!��S!��c2?��>�������)S?2E.�s`�>��>N]�;S��>�Ѧ��SȽ��򾿺{���^=F}��P�F�Ɵ�8ׁ�[�1�=$��k̾�,ƾ2�?(w�>A�?��?���>��j=���>�c��u�ɼ#�ȾN��:?��K>mp@�[�Y>�
=8 >U䣽 o��cL��\�>���X�K�"�?�٘?6�
��i߾Clc?rsؾ|Kd�]{��4{�MS<CK���Zm?�����>������`>
��=J�>�	����d�

 ?��<��=�0?�5�?�W3��Mi>�Cu?qOb>j9a>k�?�u�?��4���>ӱ�>��l?��+��j ?��d�!�(�#�-=�
?|��>.҈?��ܽЕa�M�?X�D?����^.�%��>G"A>Ҭ�>��#�VB�>��-?uZ?��q�k=�>�c�?�0H��ݶ�`�>�D�?������"���>/:?f����8��w�D��1�ly�}�ž晛��V��>�>�?�9<��@3����>!̈́>�J9�+����߾�lU>�����־�%��	�.о�^��R�Ҿ�!���ǰ=ԁ?K�>���L���<>-��>o��� ��(�>���[^��=�>��?�2���>�l�>h��?����ǿ<O ?��A?כ׾l$>�'�=�h�>r\��YM.��<?A�Ͻ ���d��é�> t%>w>,?�����"�>B˽kLg?Xi�>ۄ$>LP?�U۵>���j��$�����g<Ev*?�ia�6qS�n�!>�x>/���`�"�g�㾶F(?:�v�E���<�e����$�t₿Y�� �J?.Q,������F�=ո?H�@��ɾO�t��>c"�b���}|ʾ#'���&�=>�>Q��?�����=l�Ӿ�o�>_�<�PF�A���G�ӽ{3ξ(M�>9��Ƽm���%�4��}lV�<�>񊑾z�C���r��M�>a�,=���_������<�>�#����=B�+�q��?^�=8�'��ذ>�y,?)�侵�Ǿ�A�%|>��.?�?D%=Ǿ�!>0�۾��Q��;U?��>X����3���?�=�4�k��w,=F�?�p����>����D?=�k= b�J��8�$�����˿�u=�*���逿sWT�:�6����C'���V�'Q��d�>����/�k�U�QM�����r�����S^?;VP>�r�?���=��2?F㔾��=e�X?\�?�B��������>��3�c�?��=�Zl�����Z�=�?�0�=�	���K;=s������.Э�=�?f���2h����>/��>����>V"�> ���8�l ��Ƒ?X $�7��_�T��Nv>Bj`�A*���Y��������>��I��<�>�$?�?#��=vWI?�?E?%�R>l؉>hn��d�?�(�b�<<(>?o��?UZݽ����~u>�=F,>�6��^>撐>T̄��}ֽa���X�X|��`�t��>	>Yپ�g?��=Y(�c�<��鎾�<+�Ľ��=Y��>��B>?���|b��{�>���p�>���Ȳ<R���h�R����=�
>�����Ƃ��ʼx��3v�ӷ����=q7����/>�ƪ>ݟ2���e?i���K���4�����<����6W�=᧖=��
>o[K�b��N�>:[b<��=Zc�>�i�P��=e�=��G>�5B��RH>��>�͒�|Y�h���+�A��_A��0e�>��Ӿi�&�8�w=�*P?�3�������m�1�?�����r������>G�>��)��I�>#?�)��Ж漴f�>���>�O�4�b���㾁F >�ƾ��;���=��/>�c>�/�6qq������p����r>?VD����=�-ͼW_>O.���5>�ٿ��B�����=7f9�ِ��f�>usm���?��������w�>=�>̰��k2��j���6�>ԕ�����������>ف��)ľ�Ӟ=�u����>(nt��>Ҿ��@>V->��F>��=H(?i�>�(<�b�ž��Խ��ʾ����b�����7���!�x�>�=ǼP������Mh��Բ">��f�cJ=ȓ>��?>��=��^��>��=��n>��(>C�I?O������=-�!�Z5��t����
8>��6>:gb��FG=���>hX�<t���ؘ��?]xɽ����?~(�q�D>ƭ>����S��O��>M��=��>/$>���>�<�];���=�R���"nz�Ð��G�Ծn�>p�'�@&��(�g>�4*=��d�J��=��O��λ�,�-J�>��5�f���"���>�<ּ�d'?:C��"��>�Ħ>�C�[p�������>�Ą�÷�}����|4>J��&���7��=���3P?���� �#=���>�u>b��䨚���>�6�;2�>��<�t?6(�p��>cs�<�<_�}_ھ��>���=P���}ce���S>�L�%�'>��b��Sپ��)��M_~?x��н�Q�<w�>�~�j��%�>�G>�A����>#�;���5>��= �)=4��>�/���mM>8��>E��>0ɲ�;�h��m�>�P�'I��[���<��<�W��$�ս+ł>)H>c�A�x>n��>Xy�>>h��N�y>*�>����Ȣܾ��q�B���X1>`�پ=�<����ھ]��>�`콌*P�t�L��-�>�Ž����?�f=��?�*=Qj�>a�>���>��&�t*�QK߽�9�{��>��!?��y�љ!?HM�>�x>��=B��׈�=Lk�=�W��"�^����>G*�>��S���1�P�?Srt>T�>Vxƾ�e;>��=�y6>�I���ҽ�Q�>�^�<XQȾ�{%�¦>ԥ�����>:?U2��d��?��?��<�^	>�Ҙ�o����z>NN>˦׽s��<"�=>˘�>�L��#P>rq�?�@��}x��E�=�<>W4#>E���}���j�o����>
��=i�K��Yy>@p�>�C�e_���?x�@=��\=\.1���n>���4f�;9~��:��=tN>�׏��|=]�j��5ѾZ��>"_P=[���L���==X�
���=$˲=��d>ȷ|<��2�I��>�	V>�{���J<#4x��"�>�Bu=3*>8���|/>�m&������2��a���6l��ż�^�����l�@�f�H>ok��&\=��
?O�)>ek>�+��N=�8^=�\�I/��d�A>t�>�ʾdfP��ś�iҦ=^� ?}_�;�]>{�<��_h>��V��}��֠>H�)=R��� =���p0��%�T�,�*�]�/��~w>F�>|��>6�<�8>g�b>����h�J�>o�L=�\�=<�e��7-�#�ɾ�=�>��r�΋�=t)�>��=��=㛥=��=�� ��e?�ZK9�F�e>�V}>j�ľ���>�ֳ>��fy�?1?�[�B���>{U�[�?��bý�䀾��>�?�G���W1�P��=��[?�`��b�=��>&?�F���r:5/L���G>��þ���.}>�D=
G�=)���f>yqo����=�!L=]�����`<���=��+����>%NL>�=�6=߁E���0���������x��;L�0>L��<�B�>�K2��ٽX�]�>��Q=;s]�pg��!N�>�)	��bJ�n�E=9_o>��>���R���qw�>Z�׽���5~�/��U>O�r >�i<>�BR>�|��� i����>��]�>��>�w��>����1	��4��𵾢c�>��=��k>L���F*,���>��>eLf�3J>p��۴>G�=�@d�=>���<W�l��S�t��="��d�勼��i��ғ��r�>�Z>��ý�P�0�>,�d>���>�j��Z�><�`>P�?������!=Pn�>���;��9��T޼ӏ��B�i��;�5�=J����>���<�����3>YS�<pW��V�={��z=��}㩼Ò�<�J���?Ne8�!�e����S�>	�e��?�-3�sT�>�s�=�u��qSl=�>�>��e�գ,���7�mt�>��|��y��qN����>
�z=���B�<Z��>�i�>��>+E>���>A̭>� Q?��=���?� �r����]�>�
7��
����ϒ*��ѽ�?[^����y��=�b��>hA��OK���U���6>>�k�%��>*|'�?μ����!���$l>�J�ì��-2���0�Y�H��>AY/��eG>Px���nV>�S>���=`�]r;��3���b�A=�=*O��rl�<���>-3��-1�'Y>�S����>g��	{y>V��=���� �s�Z�inz�r��u�=�v�4�_8�>��>����R�.��>*��=Q���󄾄S>� ��'��]��a'z>�3>a���#�����<i�>?<(���U�_�=�%=�YD=O��i�>� ���һ�5��=@E���>��~��S>g����t̾[X>kBo>n��zu#�-f�� f>�\�@NU��H<�ȣ>�K���,��щ7>+Ԑ�@����ɗ>����kO���?x�G�>)69>���=�����`��g�+�=<і>�f���,=�W9'�?����c�C�f��>Ďd>�Y=�����>� >=�L��Aqn>�=�>V�ƾ�7��<a�>S��<Y�(�n~H��7%?%��>,�>$��c�>?��=�<�p���q����}��	���>����龣	3>s�S>���c��6�D��`'>�[.��� =B��ڜ�>�wA�>N�1�`>�w�>Z �={�;�S>� �>q�����du��q�>�%�fw��e	����>pKϾ�f�ՇZ=�`��@]�>}�H��1�?�^���9��:x=��?[�����,>�P�>~i4���>ڼk>�煾B/>f>J%��u����b>[��=G`!�����W��:P{y=�ھ�_���x/> Y�>��>.��=�>��>\e�>�k���??�Y>_� �ɔ�>�k(��L�=!���N���]>(��=�,L�-��<\����S?�4��9偾$8�Z�?�l��{
�8���uR�>
�G�f.�*w����;<����ɾ�򏽞�?�Z��5۾[�<2��>/�پ��M��MʾOx�>UԖ��	;��>�;u�>�`�#�ǾV/,;yɵ�a<���$�Ԑ��;�>�n>�:"�TU�>.�?FR�=N੽G5�~%�>��>���=FZ�x�=8�P?K��u;�?$#վ�=\JB=R��>�d�I )�o�j>s%2�j�G>t�=�M��2>�i�k�ξ���B�=�'�>�T����Pk����V
Y�����޽tc9>r���T*>�/s��H?�v�>*��>p��>*.ʽv�$?i�?�I<>`�?S>�L�?q��>�r�>�1>��S?y=�?E��>�q?��=X�??Sj?��>��>.a�<���?��>�l��<��2=5ɾ�_�=�wg��ű�j�
����=��}:*x�>�>rU����?(}���lN��&�7��-?x��?I��3�?Q?�����=��\TG�`9&����u��>���-�<�<Ѿ�T?�t�� T>��=~5?'���²>]�l>+̌>O�=J*��>���>�9��'��r	�>�l.?��T? �����9?GR�?ig�?nM��^��vkS���Ծ���>^HM���jZ=��N?�6�>d�M�����d�=�X��?��:��?>��^4	?��<����>r/w�dS��٭R��ɾ�Yܾ�(>-8>��j?E��<u�M�=k>«?��k�|=.w���` ?��5���=�;�sg*? w�����>j�ܾ��?���<rK�%Ƹ>�D��e뼙��b�h��<M��=�z�����h�V%>�Z�5'�j0��OQ}�ؒo�{���d������0��0�/���7��v	g��������$����ܾ ��<-4�?f᩿9�����
辿m�??���$5>B���y�>X?>{y��Ę��7��=:�M�6�ު���K"�Vђ>>ng�*�־�C����&��XI��;l>��=�V�O>�?���#>��l��=����[��>��8�U>���=����^��=�F/��ȿ>��,?�F�O]���>i�&��Փ>�"���_!��������+�"�d�� �˖�=�8"���=>�׾pُ=z)?>����"=��H0�=�>��>ۋh>�>�>\PK>1ن���>\C���/�E��?�ރ�q�K���E��� ��z�Ӟ����k>�G�<ב�l�;�S?*:���#?:ű���~�� ����i>��> ��>�4����#?{5�=!�Q�R��?l�?�X�=�(��:����,�]dʾ�.��1IR�F����w���g>��?�龓ܾ�p(�&�>�&j�-}�oF?gV~?�G�>��>��<�+>+����{����2=��>Y���{��`$0��a�	��>Gr���~�>�@���C��r:�Eҭ�VD�=��<�+k?"��>X�!�{�.?�����>�>I�(�>�%?��?a�L��>�Ъ>_�u���}����<Ý��:O?�;^�jz���>�劾G0>��y����>Z�><�x>�¦��j��H�?���˔=A6�`Ы<Jھ`��`����\��d"�X�+��(�>�����jm>�nܽ|���g������N�>�����G��ʯ�>�Y?Ɓ�=����]�?>��?��	?4��`=�7�Λ|���>?�r�>>��:|?9ľ�ݐ?$�����=�8?�#)��>�>dt����)����=?�Mؾ��?�(N�`g2�oR?ᖮ?C��>vr�����Z?�� ?�-><�?	\���	�����zA���3?��j?+W>���>t�>��m?�l�>yӀ>jF�=�=Q>���>�K@?I�V=2��=�^y������ +?\ �Kz��1��?�cؾ��>���+���8u�>�KJ����?�꿾ap�>9�?�.V?������?q�P�&��=��h?g��?���>��~=�~�>�%@��>N?U,�=	���="��z(�����c�E��>�Z=���>�ɔ�8w�������=D�_��l��Ͼ�\�>`/[?_�׾6t�����"^�>�w�s����M�=Y.Ⱦ;$=s'E��(��`�4�l6���F��	dl>G��T�n�4���?4
�&|�=�� �5����xK�S�<���	>�ߧ������?dM��SA*����4o%�3��>|1E?t��>^�:�$�?���3>=�7>��"?���({i��Ӿ{�`��Zپ)�Q�+��>�mW�)b�����%?�����,o�wk0�E�G��\�����>$5�3=>��<�/?�+�T�?_;������_��&cP�[i�=秣�2о}s�>�v8=}Ҿ��@�
݄��,_>�#�ԃ�3��?��1?���f���ha�5��@)Q�Z��M'">*%��O�T>o�ﾅ���=��.>����+?^��=`�`?�˜�$�>
���s�; mq=�d?��_�h���ێL��C?��+>���ξW����Ⱦ9~�ԕ̽�����u�>h�3��m����$���嫏>���y����Ȼ��Vʾ`���ȥ>�T\�؛=��V=S�̽M�>�����O��6?�[[��o�>�����.��V��}G>Z��><폿�0����zn�>��o>��C�h�=��c=�L߼����H��<�k>#�i?G��"k"?p��g������?-:/=�j'��>:���? �V�g�%?.�Z?�z��0S>�]�6�_�=m	���<?������>����k~��e��>ۑ>1���+F?�`���>}ɾ��M��j?�z��e�?<?�:?��<��+?���y��?+�|<��q>5'ÿ�)�?�$?ҋB�7�l�j0@N�>[��>Ƣ�I��(>�[>T���������<j�>�����T9��H��?��
��&�>r��>��?H��B�S�U�?>���
�$>�r
�ˇ�=�Z�ޗ?��}�=X5�.�J=Xe׾cE�>Z�+>��k����N��Ⱦ��v�������=����M?S�1�^�S>Χ�>�
�>��?�d��>�<?��>�Wa>�1g?���>o�?�Z�d��==���_�-�e'?/����]���=�<�ݾ�O�>hGp��>�ب����̾�?=��?�������ٍv?�zH�q�>�(�m�u��ɨ�r�=�B>���
<�T�P��F?����+;?魛9;vA�&>	�]04?��>���>�$)����=�0�>�B?mc<>D�?)��;�������?�w ���>
×��;'���2?���s��>��>~˲�h ?g�?���N@?G�??��/?X��j�?��˽T��>���>�ϼ?d�>�O�>�����?��?�ֻ>[j�>�����پ��7�>8����!?�}.�"�=��1>5ɱ?���<'o���~�B�%?}4Ӿ:��=1�V;�x#��P��%���1y>p���2�\>��=� �����c��Y^�=}�=d���á����ykξ��>'�����J��>�=�R��g&q�C�y"^?7���&�E�O�y�Q��>P��>�]I��_�1]�>�SI>�d�<]껽�����>q!>���-*�?g�=#$D��t?��,>ʦ:>���*])?7rL?�����hF?�&�yV?D���~>�Tƿ�?E'���&��#\�.`��)�J>|#%���M?�MC��� ��.X���;ǿ�,!>#ܵ��@A��񠱾�]ͽɐ��9�'Cھ����־)�0�n�����	��Q�>�����$>S��y���%����پ1��kr<�~�Ŀ8��Jq�>��9�X��C���Ɂ�Xg���G�5�F?t�w����>��U>����X�
?i'����>Zg?�2�>�ѿbc�������L���b��K�<�ߪ>���?�^��1k��]B����<��y����~�> T??�&&��Uh>�D�>:�=�0��<��=� �;�s�>����D�>:�B>�뾍?�㣽��?�W?�I�=!�=Jh>?�D �ɔ\�.�l>�"�pL��$���?>�Xl��������]�_�����-��)8��\?�U��i>����>��O�����U>ӳ�>u��[���a:���j?PJ%��e�A�߽ظ9>z>7[˾�����Ȁ����>�PѾ����:=��P[>:�>ʼ������@w�>�k3=�E�>�e4?�~X�5�I?�#*?s���ɍ��/�F>2��/��3��l��>��>\�?�A>UO?��0�Q���B����>�}}��#_�j) ��f6=���1;��!ճ�z�>��?4��>,��>�~�>d�P>8p�>|�>:�>uu�>��?�h?2:?�z>Q�$?�(�>~���x�>y|?o�m? R=g>E6��ZM�Z0=!)�>V������o��*��%D,�XH�0�=�'>V@�>�l�>���>��ٳ ���<�U�>p��7D������p]�>h;޽���=��V�H8����?�I�?'@�cM�F�侓��>�lҾ�%���w�<V&>�ŗ��˽�x>�,�>�dK>�8�>�<?-�?@|�>�z�m�|>4�>���=28e��弟ަ>�:>a��=��=m�<��Ƚ��X>
�'?@ �>3�����>�.н�4���	�z��>
��<�M����ꌖ=cg:�U.���>�#0�9�=Ԉ&���e�/(��b���??�̆=B78>��<>�P(?K�4>�ˣ>�f
=B�*;?���􈔾4Y�^��=�`�vn���玾ٟ�>m砽�W�=�7ɾP��>�G��'kq��D���<�s�;*.E<dX�=�U}� �h=7G������оr ���޾���A~���C��*-�7<�����=k§<��
�kQ>�|�7��R������"��!��>�>����^B�sM?�Q��"���@��m>1�)>��n?}�}?s��>���<%MK�eަ<�0����/�R�����¾Ȗɾ,+�+��<�w��2/>�>�R=>&7�>�Y�=a�ѾN���v�Of>+�o�� ��K>_��>󷌾�h6>�m>~��>�V��$�>/&�>H��>�L=⧥<6��>�>>]#�/���k��.�������= H���)>cW7�T^�Q(�c,�AQi�-����Ʃ>
p
=U@,���,�0T>e�>����/�>^�>I���	>�>5��>+�
<�b+��>{>i�;���e��I��hs��מ�>�B�>r [����G�"�@3���c������>`-�>M^�*�>1��=V��=�O�26�>� 	��o?e��f�!�c?><�
>ƣ�=�x�=�ι��?rJ��D�l��֔��S��s'����
�`#>�]��i��=�XI=���>*��=�^m>��=���� >lA�>��'?����=�n�>�7�>E��"�+=Pn�<	��\�����(�R�VGY�M��ӑ����ԖI?Ķ;��Z�2�{�٣??�Zͼ��>&�>���4]��|��޾�ϓ���=�'�>�$�,ٶ<H�?���>�ܴ��s��_ ��he��2��C�%>*�.>���>��=kI�=Q�j>,��>ޖ�m4a��o>ߓ�;����R�x����>G&�c��/�>��Ղ����{p���9���ڀ>���;,�ƾ��<T�>��>�W)>D�.?���>%�.��X��*���־WRa����=�ܒ>ۺ>��<�*x>��?)V0?_>�>-�>>�g>�Q�=h�����������>��н�>>MP�>�k�>�����=����>��
�(��>���=��>>m����6=�=�#	���q��gE<��>k]�m�&=�=̠>He-?M��>���>1�>���>p¢>�{>�@�>T(�?�蚽�@6>�i���z��O���[�L���E���]��!��4v�Z�������V����<���=�/�=�dI���L>�:|>\!�>c=��^K�>Zs�=��>8e����>��>�%�=d�	>'	D��؅��M�=�ռ�[ɾ7����`��i�X>x�����d=L?=�v�>�C���?>���=.�=�g�>4�?��ü�0�=��>�Q����%�u>�XV>2�r��D�ĭH�t�H=���wl��%��H�9�u����#������=������=�2�)���>����˼X��+�=G�<�X>�u��w���&m��$>6'r=Ǿu��>q{?i�=w���R� )�>]���I$v�;K���0>%�ƾ��*��iϾ#tȾwW���<�l�/������>��?R*ŽA'��A>R��=p|�<YB=��Ld�$�(�x���ng���=7�E~޾>�B�
w�>��ʽ�⨾׮��'e�~6����=R!>G�'`�>�����ؙ�k��>t�����>��l���:�ۼ%�վ�Z��1�� �;�oҾ6x>��=���v�	���>j�$0�=%j�=�~ ?b�#�e��:\��h
?�;�=��2��Bg���@��Q�=�3"?6>������W;k*�n���6��t��FQռ4����z��<qu�1a�<<{�CSJ>�:[={�<z/�>Qӡ>�F��^>B��>��<�%�I�hm9>��=D�̄�=((�>��T>P!4>� �>jq�>h.T>��1���{.��ܐ>�}���������dt>�p7��a= ����}�m��>M�2?'��?WႽ>8�>���<9>פD�-�/��@޾���u����5���A�����6��Dg�>_	�>by�>���X�>d�D=Q`�!�5>�
(�g�Q��]6�j%��1XԾ�93���w�j����m(=[�>~����� <���=d'?�6�x >(>�]?�H��z��>�"n>KeY>�"0����=��?$M?��c�NP���䀾ioJ����/��^ST>���>�UԾZXg�G�&���g���>��	��u��l�>��=AE�����K.�>ͽ8=G�ھ5C�C�>%�>�h����>C�>�e>Gc���L_��{žv�=*{�v�=�vA����=����i >�`�;�ֶ>��}=HTO?�ɨ>v�>�|<�O�=���<�7�>K	��,*�> �J?,C�>l�q>���>�0E>��=\�5J>vó���*>/;X=�?/%?p�� �>}OB��PE�"P���⏼d�"�4�WW�����ܾ�����td=P��P�K?��E?w/�r��$���e�?�����*:��p>��C>Zuž�����><}�=h۽���>��G?�L?OB�=�_> ���f�(���,=��>���BP������L��m��9 �����'%<kܼ��������7>�]�>���>������?�w->�Ճ>>���]t>(y�;��=��b�cH��?:��l����>��?/�[�i���kKk>�Ul> �L��'f�+>37���?��r>��=&Y�<Į=�֥>I?|�ZX`��"���>�4�rl���Ҿc��>��h��P�����ׁ�նԼs5 �S/ʾ`h����;�HJ�:о2���~a>�+]��̥��J��>�G:�m�=���|�c=\䫾��&��=�f�/>t�>R��@Ż���>\��>Ͻ�ⶾ��ٝ�i.�6��	�L�OZ'>kR�>��"?�釾�F�>��>>�!?�e���J�>zW�=��T>�s⾛ܓ>�6>��>=��>�aD�Š����.�~>�UX�y�����㲋>ug�L����bw���>��0�<l�<{��,R�>��Q=��/>8rg<��>,�������B�속>m���e�K��ۡ>��\�+�Ľ�e|��sp�}h���NE��������ڝu���]h?ب=ݒ����z<0d�>�_"�� �;Ѳ�>�j�=���>y���ެ�j�u���/>��O�E����Kξ���>�&����d��;��>k/���v�>Pe�=��?o	�>&z�>���>�B?|��>ie�<7~�>xi�>�Ś��YJ���/��#P���6�g��=��վ,�>C�{>��>�Z�=�+?\;4�Ɲ��4q�b>� `��qJ�𭋿bY	>���H����Q��`Y<hV={*v>ʳ5����>i$*��\��n��q~>��������5���>�)�����:�t�T>����(!�w`�Q�&<΀��P�B�����>*V�>�ś=��>>�M>�)r>�X%=�`�=��=2�G?�#�<�)7?2�I���5>ezt?6�=�[�� ���7�=����+ɽ��>��=�?�>B���QG�>�Kn���w>����������>��=�K���CT�N��c��=Ib�jO����t�>�L�>���<���>w��>��>+�=�>��>���>ޚ>�_?Z�=?�&=>	�>7�C>Z=�\<=���=%����ۛ=��?V>~�>~B>*�E? �>�m>��D�%?���mɾ��u�-X�>��-�v�>2m�>��>A��=�1�;�H=��C>-��t��|½t2�>�����{1�`	H�n+־^��>ei�>Z��=�ƾn5=X��v���w����<�a?k��A��
��dg��]>k��>N��>�?�P�>h�f�
S>y��>9v>��'��Ȩ<�Ef�6�?��
�徢lu�E���fNj=�9���s ?�ܪ�=_?.�f>�G >�����?���>g�/>��۾����?�a��n0��Q)>���Y���>ݰ���>�G6��a����<߀q>U�a�mN��ғ�q"�>��
����=���<���> �=����8�ٽ�^�sE羾6���款�#b>����|�?��F�l`�񎱾����c�^yӾ�+��3�-!�>��>J������Ǽ���=�Y5;1���=�3>�t��4�o=�{L�(��=$��t^�_�߽gk�Mۄ��^?IOľ��þ]ƾ�:?��8�|�+8����a�=_D=�x��>>��?������=r���K�=$�)?�\D>��-���!���d�>{���E>U�*>)1�>�d��zʽ=�=�i>�/���3þj1=V��>�_�w!�'� >��>�q>��g<�?�>H Q>і(>>Nn�>�.��f�=	O��t!>цA>�)�> ����*�;ۺ>ԯ����t>��ݾ;�����!��ٽg>��
��>Kb��-3�c�(>IC�>��B>���>a8.?"�;XϾlB�>ͩ�q[8>�6�h=+����*��5'�>��ܼ]$
>�G��	ྜྷ�^��Q1�Æ���!W=#�N��k#?9�Ҿ��<���j� >.K�;b>�	�>_D?UUP��k{=��>Zp�=�佛O��	���~�(Ѽ�(����`��'�!��Y[��b�<��?�D@��%���p%>gW�����>>s����;���==�8?�S>|#��-�>P��>���>������ܽ0}�>�X�>�����q>t^<�>#�>��������4=�X�>�R��?\����Z�]+H>(��>��$�rA>t�> �ɾ�p�=sМ���b>�v���`�>�䱾"7�>�[�<��>!u���;}&=�H>H��>��g����3�<�<þ5f>�@(���>��1>�����Ѿʤ=�z>
�=�g����)Y��#Ǿ:?Խ��b>g�:=�;>�:'�xɽ�<�����>x!�~%��a�>>��>(�c>��?�)?y�Z���=�I��H(�qo#�x����>��0�J��>��<&l(=@ޓ��!r>���>F��>~&$=���lg�=F��;j�4?�K>�!E?c{[>��z>�9��\u?:�,?>K�=h)��h4?g?A?^>ߌ�=��b�ǡ"�ܹ��,ᴾ��><ZG�=�n>�Z5�$��=HG>��>�� ?9��>y�?~z>=���.8?��>	�x?��>�g�==�F?�*d�w��=>�=l�>W�<?�%���Ҿ��X1��Ӱ����>7b�=Rh�>$���h�>'�N>��=�~��3�?I��>��нi���}�>˶1?��a>c�>�{��Z,	���<fN��پ�J���#��[�>��)��� ���_>iԜ>{{�<N9���g<V�I�{t'>��!����zY<�D�>-�U�-���Z3�<�>��>)��=����@�>`t����#�۾�0d�6wѾ�%���ξi�<�j�zd��p6��ד>��f>�D.��眽��?s9?ZF>4�v>�f=�[�>��>H֔��ӹ�	�`��0�>�H�y��F�����a!t�`A��~j=�L?md��P�'�Ω�<R9�����hߎ>����Q���þ���������><�;�r>}�E��6�>���VG�SԼ����+�������c��zw��G���͐=��#=�}=\R��[�>��>@�=��|��"?%��Vx?����=����>��޾Xu�>�=�q>��,��ye<�b�>@1>9�?��g�>�?R*�>�1o�x�>�����<>-&��+��>L4�9-���r�Mb?�J>yB����=r��뽗˞�]a+�tbܾ�>ע#>���D����Q>��	?������Y�j0)�:�|�CwA�6D?��>Ȯ�>�?��s>Z�;�b�=X��>>9>����\=C>��>�b��?:���>�k�>M���n~>g�<{��=y|��d㐾B�t=_�>�Ͼ�溾+<�;��>?�B�V�P�N�<ڹ���?�r�>�x�Ys<��=�=?�<�ox���>�u���L>�������S+��-�=��t��{�>w�>b?r&3=DO�>a��>�ξ�@�=q(>�?�.�1���pY>����p��k�.�����<��?[ �=��b>j���?�鷾-��>�u?�&�>�vƾ�TM>�&?���>(��<�W#���>,x�\0i=Q���c0��羆�2�ȓ�>ӹf���>7b��� ��w�
�ľB�?SA&;6�>ne�> 5�=����O���C�>��M>����|���m>F�>�핾2����g�>���>��=��>(��=KLC?�jy��N�=<M"����>1oҾ�FO�H�	W>�k���=��>�F�>cY >��!��?қ=��?��?*�G?>��=�>h�>{a�����>��i��R��k%�=���P�>)�R>FmH>j>y�>�	�>��M��Ru>�>l�\r�>�.���50�5"���8����H�ǽ�,�K��=f)?��&)�>V�=�!�>�ӽj{޼�>?6�K?k��74�Eӛ���(>~D����=5��>޳^��0=H�>�hE���?p�[���O?��K?_�[�����B^�<��*=!�A�V����>qr=� �=e�<��`>�x0>���=XG@=�v?Et�>�y���%��"�>e�5?z�>H۾���=�,-��뽦{�Ad?TV>�%�<յ����>�>`������\�>ʐ�>��	����>=^��Ȉ�=���f{=87ƾ� �/�{�)�=͕���Ǿ1{:>��,>��"���+��ǽ����C�ӽ�s��U���&��ý��g�m���K��7���L��:`�N>�U�>f?XLa>>b�>������
=x�_d���Ͻ�>�����:.>��K�b�B?��x>SbP��N����?�4?㊠�	�w�����C�<P�>�ݾS�>��f�?)p��X��>a��>l��>�gԾ7k=�D>>�i�>p���z늽Mͤ��Z"��'���8�ĽvL^���������>���;M�!#,�|E����>7�2��%=�?��9m>�<�y"7���� p�=E���j�
�>R�>\��D��@>�T�>�y����>*�S>�4��kž8�Ӿ�E)?�`������C3v�p��l�`p
��l���~>���>F��:L]��佳bC�^ ��I<���%�}>)\c�%N�n���6��>��پB^� �7�β>�56>.�9��h�>��$=�*>�a=�P�> (�>s)�>�$�����7^?ݒ�R��>�(>_�9>'޴>]Z>��=n�A�]D>��b>��d��N�=	��mI3�8��_�%?���;���c�Ⱦg#k>���t�p>�j�v�=ӓ��cd�5���8�>F?�*Ⱦ9��6r?�n���  ��ȹ�*>i�I����ş��=ݭ�>����@�=����l����	���s<���>ĭ�>�U>T���U-���a9��I�=�\0������l
�bv@? ��$㖾��R>�@�n>��8�k�a��v�>̙�>F5"�� �>@MC�.1?�V���!����=R�"?�n�=�I<���=1��=E���&������	>��?M4��_>��~>�ȫ?��?^n?k2">pA�>�@?�qX?ӱ�>�ש?!��>�+?���>L����Q�=����h/?$sr?n�>�u�?K�>�ً>�?�t��{X����z;��<�B>���="c���Q>��K��t`<��n��>�>3���R�>Z��fse��t�>���>�b)?닐��.�>Uv	�'���J�?���?��_�<�d�A�G�<'�q=◚>!$G?�W�>43��Մ>@Lc?�Q>M#���F?�/Q?s�>7����E����=>&K;��?_�4�}��>�_>]�?�U	?�@#>{*�=���>��!�����g>���E�>Sؕ?�P�=�7սш�=?������#�(�D�g?1>�����%��a�<�<��	b?=\xS?�)>����?z���?$�Y?�Dv��kþE�C?<T?3�>�s(��ml���g>>�����
�$��?��;V�:��h�{��>^	�=��T��a�=~+@?�S�=���>�l����>U�H�������*��]�QZ��$?��@H�������>�p��w���oj����4�3��_.>�o>�Ss��T���5��d��H������[ ?;�n<Lu>�݌��y�3?��~=�.�[ ���Y�=����l���Pn>m8�sZ?ԡP?Q�Ҿݙ<�����e�?A�(�,�t��[%��3�{ߠ��xϽ#�����>�g<>�����Eɾ���Ff�-�庠��R�b={��>NN??��C?��ž���[��?䐸>8g�>����U������V�W3��4�����>#��>�嗽׿>?��\���&p�����Å��R?&'?;xǾV�ܻ����2E>(i&�<�܈�5��>*na?�}�?�>���?�f����}��3�?+z>��%�<�M#��W0?�v�?��Z�~�¿*q���w>1��>�g��&?�gӾ|p��r��� �?ᘉ��EF>F&�?��?t���}�Ǿœ�>?�>�����!>3�n�G9_?���b�E����(>����X�
�K�>�J?�ḽ��>N��Ȯ'�m��"��(���Ԕ��^�?*�@�]�񿿿��žU3P=��T?�:���F(?#���D}?��B��!��
���Q�ǃi��qQ���<ݕ��O�?u��>����f�����>6{>�(q?��.�4�?�FZ>V0�>RR?��>�W�?��L��Z�Ɩ쾗��?���?�->>,ޕ��0q>o����X�>�.�[k�����=IZ.a�:;`?��>x[�#�>�C�,��>��L?��4����>cB罾�>�[�}�i�R���S��"e��$9>H�^���>��l?n�M�
��)���ҾHoٽ~8�=�����>��)?�&?}*?:!?��z�� V?Q������kLY����>U?�O4����:�F�!��gn;?HL����5?��=� \?I8���}�>�.>|��?����լ>���?��>�T<���>u�?��>�f�� ��>�Σ>܅">?���@�s�V��DN?��>��>���?��?�b�>z����<�iA=�?HfC?��a>;j?���M�>?:鼼k~?��=_R@�@-"?��B;���>�ʾ"+�kڼmDҽ�?�h�=X	���@�����=���>}@iO�!z =�)?���>_�n����>9c�?,E�>�"L�bB�>lUG?i�5>uP�=��=1��d��3r㾅zﾚ�L>B,�<���L�<z�5�'DB>n?#��j���Y��8>����i	������=?8��>`K�?a
�dا�&����T����=���>Y���+�]�q�������'���
�>n*�>{�Q?�
�=��U>h(��Aо=���Ծ���+��V=�'=�V�6?��վ9�i����.�A�6�b8
��X>���@��>�?'�>k���*��
�A���>z������8��&Ҿ��3?���?��>���oy�>X&R����=ўv��\1?�2?x�=d)�>��\>�]p�J�;�񭴾+H�:�G�>JU?  r�2%�����rm�>�邾���Dx�Bj�� ���1����w�\?��*��~>�Q>�k�>Sp�ిP����뫿��پt�*b��.�B?��>=nT���Z�>&���l-����?N�=Zh�I'��5��>��>�eX��/[��5?N�9����>�(���]���>�%5���Խ$B��B��d�E?)�y��0c�W��P���YWH��~��>S�=4�L�A�E�u�?���W���&x
?�1���c���f�'>}q׾p�I�񤑾
�?t罪��>�X>ŷ�?u�2>�H4>�?���0q���A���1�2����.����3�>ię>�w>G{T?��9�e�0=t�=�8����?_�w�Br��:���k��$��?d5g=��7����={Ս�$`-�⯿k���C��=�?c������O?��%.�?Y3���>��Z<zD����h=��ѵn>���>������
)(��+�?x�,@l���?>�ݲ>M�>)����>�/�?�1�>�n�W?
��>�H>
Q��p��܉F��, @-�W>�!������-U=���>�9�?�.��p"1?�Ҽ�J�[k�>M?�L���2��'�=[*J>���i�[}���Q >7<������n���?	�O=���4K>�?�w�S��>\�>(��e|��}`�8�,��Ee�M|־v�W<��~>�:�>��>�mf>#��>�3E>�Q�?��Q?�?%X�>/�??����4�m=t���m��<�ϾA�?p�(?��.>������x�,�m��>AW���H�0���{��={�H?�I?M ��& ����)��W��N+���-��`X�\�9����>��J���5?�@��վ���>ο��FJ?VTӾ	�>�?:�+?:̾�e:�Ap>����P�e2�?�P�>Eo>�]�?%^>L��?�q?�Z><��H'�)�,?V�>H��>��f<�"�>W?-4V?�:�?̑�g�>�=�>??_�þV&�>�s�?8��>Yd�F*�>�C�>��W>DŚ=���?^�5>�j�;��>"*�F:?��>�>^�u��l%?�Y�=%3�F�i>ʬ������XdϾ�� =c޿�y�>Ʊ���b�J"ʾ�4 ?Uܢ�WK����x?E��Vbg���������Z�n��(�3�^�{T��mf9?�q�>ɰ?��Y>5��_q�>Ǹl��탾.�=�>�h6O>$��n9�?pU'?���0�?�%?Z@y���3>��2?��E�ҙ�?��F���>�8h>m�Q��B^�V���?��>V��=��(�ޮ���?D�?����xa�r뒽���>�1$�P�9>{�y>5˪�D�Z�6Vg��ń��Y�qz�˰��.	���Ͼ�%Y>�Ⱦ�����۾$~�>���k��Z)������>��4?���>�>AE���UQ����(>G�ݾ�֭��㔾��/?�o�vT8��E?�|�v���c����?�s?B�>���{�w����?k������W]���?2�M�7�>����'�C��>f̣��s�'�y�ٜa>�	�]��I*�U
?r�=Sٟ��0�=d�I?� �>��b����>ڹh?I+�=G8�>�R?���?�>jL>�AP>�)e�ks>�u����>�Eg?U^�J�>$��>$K�>�q��DH��������?ĽvS�>�{�*�&?�| ?Y0~���$�z��?�`�c�!��'�iٳ�g����ܾ�-6�Ii�>_2\�N\ÿg{��(g?4M�=�YM��w��{�?hȰ��q]��-J��ϗ=y����a_����?�8X?���>4�=����`tA?�ܾ��A=J�-=�iR?�?bM�>8K�?�^�>e�?J,�"v?��+�.���Q�����=����x�=��%?�}?�J(��ʿ�����ҿly<?�^��4o��� �>�?��&��ӫ߾�AM�Q�->j>��	�M`�j􈾎 �Ib��	{S�B�?�˰>T�>_��>�H�?lG�>w�R?t��>~��?H�	?�1e>��?p��?�Dq>�C�<���?�a]?i��>c?�!@?��w�V�>���\H�>N\9?@6A?��>�F�>�r3��t�;��Y=S%ZI���2�'��[F?f����(��z���޽�RB?l?�n���+?Z�+?c2I=jH]�t��>�ڼ�����Br�w�b?��O>��X�M94�y�	;9�a>~R0=3f����=h��r�!��	�&DN?�/�>�*>?t�>�A#?�a�=y7|�9]�&�>	.�?9��>Or1��>;��?�]�>�3��$�Y?��Ծ�ŉ>Th>+{{>^��e}��(�>����C�k>��>��f?|3�h`���+�8Ȑ�CM��x?6�C�o/�qj��������>�#��lP�>�ľ�]>ץ(�G)�>��?pp��a�=�W���R������d�	�S>-.��G =TľWG �E`��@S�<�y�`0�>d��=�?�L��,�\��D� ���$��Ⱦ���>�Ț>��8��������y̾J����� L������o�??]�L5)�sM�� /������5��~,�?U�B	���þ����!Ԧ�M�X��J�=*�ƾ��K>)-�>�񀾀�0��2?�!&^?�a�=(F�Y�p>˱3>dZ?8[A�<���|D�Ƌm�\�}��-Z>�����u>��>�?0q���ɽ3�l���>�䦾�v�����?s�>��V>f��3.�>d+�>���8i�>�r?���`��{����$���`��w:���=�l?�菉 �/=�i>}?����>8X��N �!\B?��:?�JA�����_?����4R�^�Y#)?׼�>F1?���>�.?Nr�=����tg^=0�&>Nþdg��DѾ3�e>׷�?%�]���;
r��>K�=b4��/���:���ZN?fu�)�Q>b��=��w�QC�;LJ?�6�>�?�>=E��>+<}����@�۾nI�}�8��Z���� ���;=��ѼT@���4��?��v��n�>�����8��3�A���Ͼ�@�>��I��?�o?�Vݾ$P��!K*?�J?�@���+½F��>��?/s���PH>�X?�?1R���	�>��kJz�25>�0�>x�U�E�γ�?�����5A�Lh�>_h[>O�>G���<� ?���>��r?�X�=��о�p��Cȳ?6C�>�ړ>�uD=��>@ �?������-?򪮽L5��{�����>_K�?�!>�uľ���>T�R?�U<{���+���'?F�9?~J��<^P�Ry���Ҿv텿���>L��xa�
�>)�?l�I��Oe��6?y��ռj����,�>�?b?,��>ℾ���?HW�v*?�|������e9?\��>$�>��0>��D>�@|�a��<�[�?��>�SJ���<�v?*E;���?�>?�E-?ɝ>�#�=�5�>��*>a�0?ܿ>��=w��=���<��f>���=`>/I���N?Mh�����>f>�W?�Dt?�hr?H`�>�fS<���>�՜?���u��>�u��L2?Sb���,�?Ї�=��?��"�s�J��=J?/��>��>Qi>�yK�T�?@�>/�
���r=yR?�@x�}��?��$����>��s>�G�>~c�>���=��5=
-�>�>�X��z=>9�.?�>{f*?.60?yV��?3��%����>C"�%ķ��=?W����׽�\þ���>�V�<<���p�M�I=���*��o`>��:?���=��m�ʣ���/,?���=	�c?���>X5n?��6��s>;��l�=g6�8v���>����O�u/����n?��>?b�j1�/!���7?s���| ��j=�P�>`���;��n3�kD,�����J�=j��׊�������#�C�.�&p��0�>�x�s�>-�'��ι���;>�e=��^�ո4>�@O�U7k?�!?��5>[��m���T�?Dwt�= ;6���M=X0� ?���T>������"��߈>�|?a�?`��s� ܾ�y?��K��2��J������ib��橾@��=��9?�芿�F���M�����8��F+�!A-?-Ĕ�(F�{O�>��M�������>�?����P?����[��>mn1���>�����:=Y��=�R�>�XD�op ?�	'?�?0���T:�ƾ�>�v��<־��L�ſ���,?�mԾdzG��䉿�)p>0����|<�ʃy�\r���R�W��>�W��	�����?�k?ꍅ�2X��>i�>�Q=� ̿L�"?�i2?$�?�+.��h?����lI��M�T��x�>�|�&?���3�R=4aX?Q'����F��8g?lވ����������#?KkA�Z��kgR?�E??�/������.ľ |1?�O����k��o:?k��������<.fb�tnȾ9^�>+�$>*�#��-�i]��'��?)��K��>Q�k=@��>5=?��=-�%��R]��M��(��>+��?1�l>��?��GY�>Ɔ�>CFA>��'=��h>���=J�}>���H\�>�U)=�7?��!�V�.��>?�w�J4Ͽ�y��8�>�ss>�j{���־|��>�/��`��Nƒ��f�>��>T ���>N  >�Ӝ?�$e��5W��_�=˯=�mK�Ƴ���@k?FK�>�V?��u���
?A��>u�!��V�U�{����>��}N�������O����l	�[M�=�&���%?��V?��?��R?@ʡ?J(�>�X5=>K?vKW�j>�n���|e>�U?*n�ʿ0�?>�?׀�>�x�>nFO�.��C���B3?Ծ�!��f�ͽ�&j?4U���>�N?}A�>pCN���Z�M�L�e�>����w�5>�C�>�E�jlp?�t��ww���ƾ@T�>��@�/;�>��#���>9t��ր�bu4���b?�I�>?=�>~G?Zn�?�x�����>A�->w?�W?3�:=AM�?��0�ЬW>0���9�=/)�����Ι�?����-=��>� C?�߈>9�~�y�����>(�I>Ѓ���=n*?�?*��>r	,����>�d��f���-��T?��d?S���ݺ�Ix���J4?c�w�6�=�L���H>G^�=�eX>��>VZ��/�=��˾^��)þ\!+=�p=8�*�S�J�Z>�7x=��1�Ԃ���ؽ��N��u��K����;��I>��??���>e/�>H�N�i�ؾ�N?���=�9o���;���<A�����ʾG-R?���>8��%�8���a?*ٺ?�#���Q�=�� kZ?�@پeU�N!�.�9?u��>���?V�?�O���>;&r���?�<����>�X���!?<��>��>~�E�z(���W��n�>��,?�PԿ,��_V��A���g�v�徒j0��������V��.=^��<��'����{���>���F斾�]_�յ۾UY��7��ے]>�S,�~�=���ye�=X����e�����Ѿ$g�> ���'˿!~>P^���_���xd�%��?@+X>J�ƾ���J'�M6��v�߾��0� e1?�d�z'��k��\4
��b?����F,�7}>ƒ�����,y��>aG�>�y-�LW{=]���>�?���>��=?�#�>�\�>����K3/>bĒ>�o�>��?Q>�Ʃ���?o?�,?�澧�`?E?B��>�&�>D꒼�O0�:�
?U%��g�>񀻾;�= ĕ���O=�	�H+�"%�y/_>��y�F��]�K~;�p�ςپK���W���k��<�/��+�R����@����L&��?��𯿾�E?��g>��	? [�>
�A�� �7_6�i�>;�>?
��(�=1A�@�۾_��j��>!�s?��$�)���o>�>w�I��I�P�>ή??�t���p�8h���>�E�ğ>�g�>�>B�>����=E�-��5.�����tZ>�r��>���[���?@=s��=�|l�u�����X���7=�:���[��?�>��R�a�>1lO?�t>
�(?�e>4�a=6���PB?� �>h >ڃ&=�z�=� ?�[�:�V��}Ὣ��>و^>�v�<x���@�j>��!���7���	���k���'>d��>M<�>T~�>4�T�Ҵ5�z� ��r=��>������~ӽ�d<0۟=��,�nM���w=�)>=��> i?�����Z���
>cD?���E�-�4��>�}�;�$1��'�tw�>�g>�D�>��?b?�� �=�=S�B���>������(S�;��>��ľ��J�ew�<��q���d�����>bqg�`R˾�C����>FS�<:����,�i���瑾�8�u��!�������)G>�X���5ɾmFѾ��>7M��9�sy"�L�B?�k�>�0��ԯ����k>��h?��?�����e�>F�;�����C�>\��>2�C�S���r�>��>�V>m��_�O����>��½�)6=i�L=���=R�*�����m"���b(���5=���>�ب��Tz���M>R&��|��Mk>;���o�=�˜>{$���g�>�ћ����>�V&�*�u������>;n��������F�>a�=>*K5>����	S�=��>{��q������H��� �>o�>�ӷ���='��=�s<�������LOپ�_F���>�x�=�J`>Ӧ�>6sE=��~�0�¾:`>�V=�|��s������=듙=��=TQ�=H9�<��>��g>%��=qѹ>�M�= 﫽�o�1�=n':�0��4��=�/�=��>D�u=-�C���&>9V>�ω��Խ�?�a�>v��� a��*{i=~�>t#̽�䓾��>h�>��=>iG]>gq�>��d>���=��r>8�羢f�� ���"e=j-Ծ�(�>�j��ŒӾ��\����˦����<����X��Ơ>&`�����=Bʾ����(�>�l'?��YS�=�r�>���>%W���2�1���/z�>%���S>}D��v�5<�f��q~���H�>�R�=�{=�p��n��6�=6�>)n���*�<���>M�E�(t>���;ŷӾ�'+>�\$�E�=���ob=>�{�>q��=��Ǿ&ٞ=������F�Sޱ�#�>�W���y��+�=}��;��-�k���P�<�;�̥���Q7>&��>��i�·�>B�g>2N�>�P��VT�/�5�HB��^:�=Tun>Ė=*9�V��=��c>3�>������f�U��X(�;�<���̼D� >!�~�m���_�2�`�>�?)|><!��0Z>1��=�����������_n�ܢS��u>����c+��L�>y%�>F<�AȾK������=�C>��H�br>���>���>w�>K?Oߢ��2����,�ƾ<��=>>H�=u�'�#8�=��?O9>�L�=,�~��~�=��>-��>]N��� �I���`l�>�����!>�>?���>��(��H��#�>Eλ>{˟���O�̄�|r�>��ƽ�>o�����7>��`=T��=�cJ?nw��]?	��=`��=�¦=�?^=�>���>���>>H?�]F�� �>�� ��e��g<�>��H>������Y>�Z׻�mc=�}�<%�ھ�o��*�ڽDx��A��=�1��P���^�>�;N?����⫾e<<l�b>^|<>S����9�[�$>�=��y>�T&���>��(>���>�Ì��M�B��=�;�>��
�v`�|��<p(�>.�3>��Լi�Ϥ޻�"U��ܦ>��O��祽ƿ>���>^�D��ƴ>eӽD�
�U�⾙��=!R ��~��fSؾ}���0T5��D�L��.�<>��=�j
>w8��|�>n�>I�@>%kK���:>Q=�>�X�=��=�e���=W]>�2%>���]W="w7?�� �Xi�aP�>��U>r4��?�V�q4<��o>-S��UC���1��Ҿב|=�S���QK��,�?��1=+Ft��k|���>HV�=�8k>Eß�9Ue�����@���!����=h�?=O֏>��ɾfW>�4�>޽)��GC�>�4��%z=��6>��;ܑ����>�V?m�Ľȵ�=4w->�瀿�c�=!_��@�=��q�$C�@���<�g�����&�c>Hs��P��>��C����>�i>��,�+��6�>�琽o���������>n>%={@>:¾�>T!�=4�Y=���ǣ��b>��=�6M�����T��=�龙'��C���)�-�T��%��ܻU>�m�>��=Z�?C�>��R�p�?�P��6���rý:	b>s�s>.��=k� �Q��>��w>a�>@��>Q@�=c���ӄ�9���$һ	e������y����h劽��=n~=�½���M>�E>~E�>7V��.���7���e?*Ow>��.���Oh�>���<���Hr_��y�lLʾ�z$��vW>�?l���Y����%>8ݘ>���>�>Z�A��"���1��������~课���C�r�|
�>���X(>)�?l��>�<ﾄv�=�x�>��
?�侇�	�#ͮ<8O�>�|�=̓/={�>�"��v�!Y����{>8���L@<�C��2̾�刾+�^��Y��J
>S�-����=���=�#<3f?���=�c�"5�;c|>t:��>;�Q��i�>m��=��>|)�J-w>���>��5>m#�l��=�2`>��}>��4�g���qA�"�����*��t�=��=!��>�G�>Q��>ſ=�%�0�1=h�M?� 5=�0<d������</�7>$��>�&�>��>�w�z�>ՈἸK�>Dԧ=�=\>�|�>Lk	<&�ݽ�G>��:>� �W8T�AUϽ[�X����BT>��.�8*�sZ���P�=ٮ">c�>qi)?6�'���>��c�>m(b?��:�xf���x�=V��>��D��0o��끾j��>z�I����N�>p}V��濾�ex:��>�~D<N!B>�+6��Y�>�+_�,�~�A=���l���ɾ�ס��?�=�D���rO@�>[??S
0�B˽5L=�!�>��S>�ۡ������=xe�=Ûo�;t�=�E޽�G9�CH���]�x�g>�6ݽ���7A�>�`�>�9j�f�~���n�u�a�H�>�J_=�K>���:ƌ>�y����X�o�<#��=`|=�x(|��E�D�'>Lq�=����s��w����,���+���3������ҽ��>��ڽ65<~zG>�� ��U��=���@,j=�=7�5���=����(�1����>�:=d49>�p�=>�x>�,�>Dȍ���>L�ҼGЯ��!t�����N�<?j;>N����	�K x>?�$?7�8?�JǾ�r���>] @>���w���"��J\�<+v�>�^ ��#>��<@ �>����|�H�x2�<�>P�C���p�W���0Ж>�K>�+������g�>�^'>|�>���<��>����=�Q�\"`�l$�=}�{�a���b���U�= >;�'��#U��.�=|�Ľt�T��>~��=��Z��t��e�>�W�=�������=��>�ܹ��K�>l_��}h>�1�>?��<b�۽�W(>���>дG�7���[����>��3��þ�Ľ���>��->��=�O�=�G?<�Y>b�">X'? �>N)>����>�f>�ᨽ�w>B��=��>���=���x�Vj�>| +>�ɮ>bZ5�>��>n�[>?��=)��=7q_���������?�:+=�֗�4����@�>�{���>�𔾩��>�9�ء(�3�h�Ɩ>Ӱ*�����!m���>��j5�ÃȾ����{���[׾Dľ_#�>���m�l�3P���>�y�>��������0>7F�>}��>x�>U �=�O�.	��if=�I�;U��>�>��-��>�Qľ�Cr�\�>m�s�1�d��C*>$�H����=�͘?L5|=�y���7�>���>�O�T7<�ߎ>`�;?q�.��;>Iף��1->b���sl��%����:H;�>l��>��>��?i޾|`о��n?B�k?��3?L>��ǽp�.?{�?��|>�|$>(�>U�?{?�Q�=/�ھ���˩�>��>|�%�y�?�e>�ɾ@]�"n�������ǽ��?O�>E9��1?`�>��K��{��ɘy>b��>��L��t>�Ș�J�/>lao><�=�
J����IH>��=�m~3<������G��_��@�����dn��6A�ظ*?Ц���}訾%C����?��V?�A����?��I!�<z�4���>�tp>S�1�vze>8�7��In>(B�;ƌ��to�#	�>f��R��>o�I���B{>e�?y9>6�8�g�?˵�!�������DE�P���F��G�>x�+�������>@�C?;X�i�S��;A��?;M�r\����>��9?��W>_����A�w�?�X���|��>��e?��L��FӾ��b�>���3��3�<���>9NE?n� >���5�㼀n�j��>[��A.���Tm��
?;.���ԾGsF?�n��(�:�%���-����>]���6@?��޾(�3���>�iQ?�rѾ{̌���=Z�?�'����M�3�ܲw?f9>�u�>�r}�f���Z\>�jN?�"�jm�>Ep�����>V��9�8>Q��?U��=��U�����!��=�&�����>�������g?
�=������p�>e��>36���=�>�`�>G����*gw>�O/>?� >�_�?ž��*2��H�=�c߽����i�@'Q>�ۺ�V&�=C��=��
�>X�k��=-2��ؾR�g?[��q̾,���#=S��&�c�p��<e?���>�>�n�x�y>��>ur�>v`�<3l==W;>�����.���D?/^�?o���\ >P�%B��~Ќ�1Z������2���>�p?k����t�y�=��T>�<>|`��m�6?r5>����;"޽J�̾0"���� ?	������,a�^,�2�������=�e=���r�">t�$��?�^���g)�����=��X?��9��	?�տ��2?ä�Ǧ�>(�����>ׇF?�ı>�+�Y*=�a�J�����Z�T��"��=L�x�c�>-�����=0�s�k�>Iʒ��{�) 
>��>� �=�z�>��>�&�>M:�>=m¾��<�~e��ۋ=��u>��R?��J�t�!��<?غ�>��d�ךE�d�>�˦>&�U>p|*��Q�>�uE?Ϧ���1>d�>9ƃ?�#����� ]?�U�G������[�<:ý7���V:u�V��z�70?b�>��;����T�������9 ��G�Nq6?���>���>�Z>v_�>%��S�վ9�������?Xx;?L#~��Y���� ?{�?5�;q#?V؏>�u>�G?_�&=�r�,��>H�?�Z��!���'?���?�x����H�>�H�=�)ʺe��J1R��M=�^?jRο����������<�!'<D�><�慼ęD?��@��B>��m���˽S�*�xf-��o>:b�>D�7>�?�8�>�풾o��߫���� �=�qa���.?C~Ծ3Z�>�����w��¾pkL>�C��Iz?�?VՓ�J���?ģ?5$H�����洿>�-�=f�?E�Z��1>0�X>�Q�=RZ�=Ƭ#��F��
?�v�>��t�4��RUf>�2�>+�=����@��?����).>O�=#�R>&�ž�C?�;���w1>�!Q>�%�>x�����Z>v�=v��=�q@��ާ�N%�
�9�O��mb
���b��o>��]�&�:>�B�>Į{?h�龺�P����>hڤ<^�0>�m��G��>�>��>k;>%��=7��$=Fa�Ȧ��F�꽏2¾�g6�j�)>-���;��x��>�K�>x�j=N�?��Ѿ���c �g���0?�ҽ Y�>��ԕ?��>��f��j�>u�/��=�0?3�V��U;F-y���x>�ic�j�$>7#\>q<v?�㜾�;��1?�䂾?D�>�YH�儁��>�gҺ���>_�?�h0>�Z�z����R/<F7�>��A���N>��x�:��=y��>JC>�O?��Y>�z���?BAӾ��%�ae�>2 �?�O7�4�C�����Ƿ�>y�Ⱦ�ɽl@��f1>��?�|�>2����ѹ�{D��`�>��Q����H��=�����F=�;/?hf=2>�|#�_,�y`o�.l��V��JK�C?}|;=u�:?��;e���3��
3?C[#=)�i���
�s��>&�S?�@P�`l�>i�>fA?�,��C+���m?ð>�����5n>u�?�	�as>!���ɨ�>8f><K��=b�>V/�>��?�eu?�|���؍��5ཇ�>p��=R3k�"�뼇��>��}��׾���������aM�d!H?��|��>�����S>���=l���� �;�~9>�[{>_��=U���썾�WP��#>wP�=��z��J�>+�?a�h���]=S?�kF?�.�;�iB�M\�>Ξ�>v�>������=����c��>pn=���><Ɂ��,�>�)�D�i�V��8-�C��>C�� N�=�9*?��¾$}"���������ν=��>�y�Z�n?J	�=��;>AX`���f>1�>XB�%�ʾ¤:?�P�>�pI��a>Z<c>	>���)7�1��<́?40�>�
p�W����?�X �g��>!�>n{�>$�/?k�>]\b>3�ʽb:�>��?��?���>�8>���>����e�>P�?v��=��P>�?:��>]����C<�E�>�ؾ�h���/��/���0��/<?ӵg�i0��G�^=<�I���m�xN�� ]��C�=i$���|�7�>*n�>�f/=����M�=�;9�+�>
ƾ�.���Zý��>w+���-���ݽe��̀=e�>i��>��������G��Y|�>��a=M�^>����n?�u��o����=�8��j�{��c���O?��)?����3�� �?Wv�?��r�{���X>g�>U�'?�����>�~[��c>���i���C#?��c��t�q�>]�M?pM���8� z<?�?	=]@¾�̸�����(ۥ��LϽ|�*?�~+������>A�i>�X���ĺ�>x�>��,��[=J����z>{ 4��4�7E�nkZ���Z��r�=iQT���\>���a�}��>�l;�)�?TY?��G>	������;>�!>�E��@�&�? �t�!�<�a=Qd?l=�2�<��I>!��>�!���=��G�>�<�M��%���ѿ�>�?t5��8;�A(�?]�3??��>e��C?�R?n1��!�mf>f�g=c)$?r��>�t`������>�B?����ܜ�ƁB>ƿ�=~r��Rt.�e%����>��m���лxO[�g&G??��R��N��>�̳>!b������>ʳ�>f*���<�>�\p��p��+���.�����;��l�>� �e.�>�&�1��=t�4�6i"?��=�!�Bd?f?���=�7b?�9�hЩ>�N�>s����m��ػ>��'?�t��z��$f)�4�{>�˷�-A˾^��>?�*?/���#/=����ZZ?'��>]�>��?��]��G��r�O��U����f2����>�W����>��>�R!�	L�=��?l���Mc=d�x>�w>����4�v�E=��/�Y�Q�Е�=����U*(�53���o�ȟ��7]�? 6�:�Q���>�T�>gsW�1/v��h�=�
?ճ=�z}=ɷ>���=>���������z!k�q�E�:�N<��>}e?�]��_����7�=r�,?3Y?L��н_u�1IQ<-��>�1���쵾'>�'�gü��X���?�6?���7'>������>"= _���<�s�Z�����;{A�(�����g=$/��슽����N��=)7�:�����Vf<�n=T1�< �Ƚ�����`�=괺=�^=�L	>�.�<[�<	>E�=��/<N�>T=�5z=F�>�[ܼG`߽E�U��==�>��=榒<���=k�=ﷃ=�9�F�;��=�<0��<��(�{;W����J���i�=�?��=��=�4U=�F�<�D�<��)��d��}��N����=���<�f�<B5I�"=������W������=�ý����@=�i�=x��.�U=��=z��=�-.;��
;p��<�~!>�>�c:8\>�I>�Z���6<>�@={��=��v��)�cۏ;�w">���?B&��4=��=��g=fC=���G�½��=�>1�=�@彽Tǻ��=qq�=i��1H��;��Ñ޽����B6q��G2��g�����7�;���˕������=��9�Nf0�1$�3��=a�=J\�=P�_���n=�Aڽj��{����<1�O��o��>�\�=��K��6�z���~�=�v�=ZƻJw�<K��3�=�н��3�?�!���<�;Z=`Ȧ�@l�<�r5=]E`��Q��G�ɽr�ǽƱ'�#c.��0=&��❧�~�߼�M� �ػ���w���vd�=�'��Yκ�M4����>���<���<��;jŔ�r>>�'��]��5'=v��=�(�=�/�_���ޣy=r�>�d"�>��da5�e�2�19;��P=����z
�JE�Ig�oX�;*�����;0�h<J@�����ãI��R:=�eL<�X�=����c�)z8=��p=s��=��ɽZ7��b_��?ͼ�&������=��9�"�=�n$��#=�ؐ;l# =l�<�i�=as�=�Xλ�Ʈ�����A�=�[=GE<�B��!�<�n>���;� |=�=�w�������21<�q�>��<�A�<��==�����{e���<��.�%EʽA�����{�C�)������\=��\=0
���<��[=��>����lCr=��>�n=�o �襪<�Z���a�=;�����*�Rn�x �'�Ἡqɽ��ؿ{�XO���!��H=��>R�J=};t<�.N=�;R=��=N5g=�㾼�@^���>���<[@�=o���=���=��<0\��Hy�� ��
������<�����<����>=���x�����>�>��<!:�%5ɼD�=I�=���=��=��;=�u����=�5����
��I]���=pJ�G^N�
Ϥ<K�F�j�5�>�:��� ��<�u���?�N�=R#�=��7��b��s�=j�<e�"=#�G�����X�<O/�=��?���	ý�1�k�h�=o̽fe�8=eB����g=��(�=u��<Gٽ��	���h�]P/>��*>1�='��=L���D=HiD=��Y�o�<LI<��=��Q=$��=^�o����<�w=t��=R�S=	IZ6�H�=X�/=��<������=��=Zޕ= ��[�=+�>�n�=�R@;qy>��6=23\=��)�kn=�T=[sI=�S<��<$�=ç�=���]v�<Z�z=M[�<�~�=�+�<"��<h/���@=���亼Pi=o%�Ձ�=�{�<F�=;
�=N�<��=�!�=��@=>�1=w�����=��V�H)=���=i�w=D�L<�h�=N >��X=r^{�[��=R��=G��<"�=�C�=�Z=ul�=qd*=@q����6@��b��3��:�R���)-��t?=9#��!N��y�<%��=k=��Ĭ���V��4�<�$�<�8��;=�L2>Z�:=)1���;�C>�q<NQ�Cޭ�I��M���X��Q����<�����y�)=!a������d��X�<��=��ʻ�Ҽ���<��[=���=)=�<]�9�#A='K���΅�Fe���ѼA�ݽ�V�;�X��m	<�r�6���<��R=�V�<��H��Ű�n�������⫽����6��r��W�¼��=�������ǣ�6��;��;��h<?QU�]ՠ��ܹ��])���齒���ۊ�<$�g/ݽ	�ȼ#c�=�H�Ύ�*��D�[�~@½:M����<������1=a2νk��<̇8���)DA��P��nL�����Ľ�ۮ�`�< ��<�
M�zϮ=����;e꽪P�=���������3�=l3꼚��g�z�=�ȶ�ј����2.�.���]�ݽT����<4�<5E����k�.ۻ�|+��Nѽ���-��g�ҽ^���fֽ�>�;T�>oE�=�μ=u�2<]�UԽN\t=!-�C���^����!�2���(���9��vU=-��<Rq�#gx�A�X�r}�����Z���Ⓗk湼�����]��"��==�mv�J{=��D�~��:(s�=�>=s�W=3M�����,���{��=Β���&>Ф=12�=�u���$�P���y���A>��=ts�:����>O=-se==nd�P;=G�=�i�=L�<T�½��h�ϰ�;������Y�����)=�'�=����bռ���=Un�=.�ֽD�=��<=gɗ=y��z�=$,=v�=gn�<�e��5ý�Jٽ�=<��|=z���p��n��	��@��=JW���z�!���=��?��O=0�;<���<6�>��N�2*��B�����;	�ڼ�+	�&���-=Ќ:=hL �^j��-R�=�=�ë�P����l�=�Wμ����I˽d�=n'�;�m��~��;��ݼ���=z�=`��=�> �\Cb=#j>%>� �<��=N%�=\pW=�驻.�=�À�秀�n�<�l��ja��g�<��v=䐒=t�c�D�1����<��<�i=����5�;�`Z=ίʼ���NW��K��E�=P�T�﨑=�k�=ϑ9=��=ZP7���|=�2�<Ŏ(>��ý�<��=$5>d���ޚ���w<(D>f]���K�<��=]ũ;7�x<%��;^=-Od��������=�a�=�{~=����ڬ��=�_�ؔ�����=X	=�?�=Z��zc�==H�=Fo(=mOٽ*>�i�=p�<�n��
K�<z�.=fV�=`����b��&�'�M����<h�M=�uw��ᇼc��TI�<�>��E<�@9=���<:MW=���<Q)l=����c�p�'�^X\��L���㽕ϯ��"=Ţ�+ܽ)��>\=��ҽ�}H�'���W���]������u��=1ވ����0t\<cUֽ�vT��-Ͻ�A���j��%W=��μi��U@I�4��;��}=�)=l}y=�j�;i�=+@e��.�<����RI=H�f<k�;�N=?3=A��6�Q��!=�E>1�=�A潮,�=y}=e4=����=�\�= �=���2��=�Pr�U����<I<����2�����z��P����.c;K1<����b������;�F����&�on=�~O�	W���U�A0�M�4�^
��`�����<� ѽG�f��<Dkb={�߽K�½�SD�c�6��ǿ�;�S-=���M��K��<��`=%������R��vo��?;R���:p�lQ�=�X&>n�k��5���aݽ�L0=�����݉��=\:�n�="y�b�����齇Oq=IO�j�Լ�\����=?>à=%)=W�<�=#q�=7�/=�ȱ=F��=�?�<���*�;���d���%"�6�3>��x=.��=���=�
>��<xȝ<d�I;��>�=��1b���2�;6�Ҽ�ҝ��#��c�S�����Խ����}�=�:=w�XU�����=¨����ڽʏའ]�=YP�߼9�ƽ�)��Y����k������=��=PR`<��_홼3����<VL;�K����=M�>K���[�מl=z#�=ص:=� ҼR|�X�����5=\��a�,�x#>�]!=���^�x������`R=�/��-������=�Q?�LϽ(�P�	���?ѵ�9�&��ߺ�[�q?>�Z�ⓖ=���T�>MĀ>Jvs>�S>��&?��'=le���'�ݽ��/�>�Y�2 ��HD>@���>OQԾg��G�=2Е?��>=N�?�y.>�; ?1i�׽L=Q??m�	?��o??��bZ�>��|�&����-�>�>'�n=�{s�d'ʽ�J'�W#�=4瀾%g>�!��s�1�Blg�5�n����?��=����/�Dx����C
\�?����oH=�"����u�����:��}��?3��>n��� ��>*"8?��>��?��? ��>�}��LýM�g��,+?��(��s�>Н߾�r�'�!���νJ3���U>��+���?g	?��������PG?J	?ѩ����F��p�?J.?��¾�`��΃i�g�^=�1ؾYO���hl��X�����������׾�?�̉��R >���>�?'�3����"�>H�>�C�M�C?�H+����>�.h��ǀ>ބ��y�������20>G���8��.���� ����>���� w���վ�j���?�=^���@=4�)?�7�95��j+&?�6�>��S?}�M>Ť>��ؽ�p�l:�ӵj<�F���'�>�̈>���=!��돚>I1=Eܕ>������(>{������>�)��C��>�}� �L�Es?�0?Ya=��8��~H?l��>z�w�컼�lr�=C��QW�>;9�	�)����!�Yx��<6�(V��V?7����=�P���u ?j��=:�2�[�v��w>�i"�E?hI��Qx�j!>?h������x;?d�-�j	o=�R?9I�?p�>I{E�}+D:��>O���~�2 �p�e?Th?˟�f���g?&R���[0�ŭͿN/�?+�>��l��r���dI?�<?��>s`�<!9]>�L�> �N?D1����>Y0���̾��A����>):?t&�>�%ھ��U�o� ��A��>^���8��'>#��?��<+?�������?r�=�)Y�@6J�+��>�k��S��|��vCP��{�<|H?|쾌3�=8�N��.�1�>tԌ=�����ľO%?w�o�F�=�}?ʖ�>J����x�>��?�޽���>6�[?������=>�-?S{�?-����2M>��>�?^̗� ����h=�8A>��	�
�?����i��u�> �����oʽ��k>�����9�>�O�>�!�>&�?�νl?/����^=�Nh>^tb�ͬȾ&#�>��>Y�?�RB���-�?s�5?D:�=z��IW(>:��=���?��=q�?r��?�|Y���>
�?!V?�XH�\��>��>b��>�@��\³>�}���0�����&?�	�0�ɨ�=�}?��Ja�jA�=��8?P�ʿ�󕿽�2�S?���<,?t'=D�X>�݀>�v?0��?�i�>oX�>�q̽�D��.>�1?Bľٿ����J��ړ?�d?=��O�`�y8?R���n���A�?�Y�w>!R�=a
p='�0�iS+>3��>ݷ\�[���?�w#?�r��EB$>c�R?���>ѐ?Q�>Y�?�z�#"q����@�> �ս����v���]]?�$d>ў��zue��T����<G�P��.��:m�>Fuu����;�l�>�V�>PȨ����>O���W�@?��r?�\�>e�? �?f��?�*�@Q�>N� ?�u�>#��>��>�m�>!@,>�`�>��?�;�?
��>��4��
j�.�2�j��?�̼�u��j��

L?�o3��*�������>���E��>^�H�k���0Ծ�x;�~�I{���<���>�0�>���N�T��\?�Aݽ�Z8�<���\�W��>��׾��׾#~��)y� �߾b�>��a>�F_?�Ib��C[>�j>�'?�Q��MF�>���<(n?*+h�v"N?U�F��x=���?l=Ž1�����u�V� ?�?��3sG��c���?��[?$�>�˾��>8!�>��>V�پ�G-��/?�fT�"� >Lÿ��?Y6�!�*�BjY��I���>f�?�'T��P���_�jb��_��:�?R��>	X�>pd(��}�>��>�~�>
�W<o{��l8��KJK��{ǻoS۽�Mq��V`<l+��* E�\F<���>�oY>����9�=4������rɾ��;�h{��O?�+?�!տ�g�=>�>��?z�п窇=eD?�C?d۾W��BKս�_?dsy�F���[��������o��T?㷿Y	���*ؾ��@=���a�R?��c?U�K�W񦽺26�e[��?�֡�E}b>NႺ�R����>j�����d��j���>��;�㱿�[Z?"d�/+%�vE��2�=O�>�nH� \��R?Ӣ���L=y�{:c?��>�A�ۋ��t??MBt��QB?2�m��a�y�����g?7�>��>�����L?��+�;
=�,/>�h�>P�?ƭ�D��>�~��� ���>��B}>�D�;�{=�DЊ��C��2?"-�>��ǽ� �IX?`����c�6e����?2*���9p�3$��p?�l�>���> ������?��,�>���a�T?����4�^>��e��??μ�>��>"U��㾆����6�����=+7���]��>�>R�M>u?{H��f�>�K���+��>�9N?�>�I�����.��?yO��н��d��xW�?$k���<�>�V|k?5$H�x0T��c�OG�=$\�A�n�W0�;A>Af��1��׾�&?�#7���FK���?��?�_X?���>f	�>�˙��N�l3?�z�> ,��+U?{1m?%���|w1�����=E�HW%��f�����pן�HP��>Y��>�ι��l�%Gi?�G>�HD�Xb=o�u?��,>@oѾ`Cq�0���� ����<S?��?�E?�ت>a�>�3�>9�����5=�Y�>�$"?FW��<�n?8\�z�(>��>�?C��=(�>�NW?�z%�Lu��;?��P>� ��(���B?�h�?�4�w�7�^&�>�)����>�?C�T? М?c��2�0>k�=?z'?A��>H4?ԧ�>Rt>���>[o�?e�g=�#k>��9?��˾s�>]��>P�9��� ��%H?㖖?a��4h��>%#5>r�>���>��]?_��?��R?)�I5��J�:n?���Yɽ	������=���t���t�d?�+��H�Y>Hab�ş��g��>�1�>@�%=.BZ?��-?�=F�g�/�X�H$�jl?g��>�Ҵ;�V��x �?��뾓� �$�߾>i�=�ӟ>_My��1����>.X�?\˶��7�=� �>ޓU?}]���B?�K?�Zm?�-���r�>�tc?Ʊ}>��.?���?�"�>0��=S��>7�Q>Z��>?�T��,�>6B�J�
>Rl�=ۻ=_N��o����K�X>��־a�����_�ƾ�eB��š�i�V�����L���iP=8Y�����N�׾���\ai��C?Ү�5���M�\��54?����^��>wK:�Xb�>�[u����q�����>���>��پ�b����?ւ�Y�ľ�1�]�?K�
�(�ھ�g�g͏>*����J��Á�*?�an�`{�T0߾.|J>�Ic��|'���l܃<�{��?� �m��ȥ}�D���q0�WDT����-��?����3;��yS?S}��j3�ɶ�>��>w�~>�ɦ�\�?�������?�%Ͽ�Э����#MR>�9?}HS?g��?�P?�ѿ��\�ʝ;��?�������:�?�o��l��&��_���:⾘�ֽ�-���B]=t��	F�5'O�f���潂D7?�Yj�F^��;`=��������E��;5L,��#J?@|�?��$ML��uU�z5>"q���H� ��>��߾v^!>�s��^N_��	���.���?��¿��?���=
x���&b�%?�ߑ�E���>i�X?�S��k�H?�TG>�(��U���Wr�>z�=�)V=bA�>�>��~>"�{�t���-���$>�ڞ�(���x��� ������ɾ�	B>
i�=�;�<x��=J?Mޒ�4Ι=e+�=�>�_>�1�o��%?�B0�z~F���q=j#>b�>�?ֺ&?��=Gjy�Au�EĪ=���)U����l�z���BHf=�sw��|��-0�>\u�<!j������~ړ>�ĵ>g^L=ԯ��o�%=yy:>�߽[�����=7I"�g.h�Q>�?�	#��y>�
�=c�G?��X�	�>�p��\=
 q�!����=��+?>.�=��(>2�>�(�>ڍ=�U	��l�<L0?;D�=|*��ʾ�j�>k�>��6J=:Ͼ��H�&�О����k�4��"1#>*��>�D*?�o�hǒ��O��Q>[�&�c�����@JM>r���El>�\w�Z�&�>� ���~>�R�����J�&�#�E>F����ν:x�����>L!�>Cxq>:P��Ц?2`�#F�h0��~�>���ڐf�_����>\;�=���8}����>@;'>A�G��{�����>+	�����`���=Z�=��>x>?�׽���_>��
?�Q��V.Q��t½��2�O�=��5�;	7? ��D�q	��1�A>:���ó�wZ��e�>�7���P�A����Z�>�K��ㆾ�þV�q=�����C=���<,wO>��>�>��E�5�"��U	>i"��ܾˬܾ�^쾂 I��}��D�����;慾��>P�= m�~��
�=��L>rH=(�5�k�>>�l@>���"�V2�>)ʹ>��>.��={(�>5QY��'�\/ƾz��>����e>�~.��d>i���v�R>�˽֡#�����},�>��=�/�>%���8��ZԾ�o��3��>�O>����k+?��K>9p>Lo�����>2�K��/���13<��j� �>�?r��=h���>v��L�4���J� 1T�����=��ھ��r��T>�MS>���=y�޾I��>�Ҝ>f�U?9�?����=>1U�>�b��wV��h>p.*?ٖ���Ծ���<�?�=����>��K=��t>q��4�>r��}�Ⱦx��w�3Z=�W�?F��>:�>];�?�群l)�H�>��>��R���I>M��>d�>4�]�@�=��ŸF>_]�a��=��<�� >�p>T�>gI?�����ٽ>�AD�+��Q��|�?���M�y>�{B�S��=�H�vAL>�(���M�|��c>O-�>�F���m=��Z����>��Ž`T�Fi�=�W6:v}/��������/�=��L�ѡ�=��|>���=ߵ&������q���7?I�վ;,ݾB��I*�>"����<��Ƚ>�錾ws>�?��'A�������� <��>腽=��c�U?v��>�D�>Lk��k�>�oϽS�=�m�<Aܾ�f���>�@�=&e�:��;�z�<�j>=�>�>> �>��=�Wu�657�(>��?�=6]n���>�;J��>=F7�y��>�,�>O�>�]�y��dr�>r��>ޟO�֓�t���0�˾�뒾��>VZ���>F���+�J>�d�>�U>/�V>��R�V�<�t�?փ��VϾ*�>*�>�=��}>�2>aY?�G����>��>����������r�;ڶ�E3>H�C��s;>��??��=l����ͭ=y�>;�E>c$x;?�=��>O՛��i��X+e>�c�>\�(<���=�ă<��}�=;��؈%��i��>�ͽלQ>����־}wc>���>惙�7�Т�>�Ti�b@0�����̓�3A>��?a�)?����<���>|=O]����ϽZg�=�a>!�׾�&�k���Ľ]t�v���Jo��D�=T���W��eؽ�?�M�<�]�;̆+>�
?�w>�[7?��>֪�>s�>rJB���<�)v���K�>+��5�#<�����w�>�4�b��S�?�rT���;3��ꉧ�T�>���>���=68+�s�����=
ع>\����3>=W�=��?磋��/��\o<����z�y��&>=�-��~�Қ<�����7�?Eľh��*	۽$��>��v>���<tP�>���>T��>W#?�F�nU!=��&=G-��o)����`S�>�i���j?��U>�o��6�Z?���($��K����c>�c��Uv���4��X�>�4
��a����b�>`��>�p<'�y��7���׾b>�����[7?c �>��>R�彲��=�Ƀ�����l񾵉��.�9�Z�0�����>-o�>��;=j�l>03�|䖾j�"��+�>ܑ>3��=%M���>@��=|~a��5���>�!'>�����-���>�R#>�mE�A�"���(>���>*�(�5��B�껚`D>)a�������q>�Tc�e�ѽ[I�=�֬>�A��`���P>V��>�!�=`M
�j�;�B����Wb�����t���� -�=�FV�hp����oH?�q%?꨾f�+=��?Ts��ʚ����N���D�-b��&H��C�>�vC?���>k�ž{QX>NM
>O5�>�����>�:{>�?�����/�� >T�>��H�h�gP�=�8�<��>ӎ�>��>�e���D=Ѿ�6��U���j�@�d��eb>ۜu��ɽ�9�>˂E>��>�x��z����|�k�>��=������5$?��R<�A������>��>��>�t#>�Z>c?&C�/���F�[�>�<�#� �>��>LӦ>&�]�F�~>��>}��>�rL>S]�>_E��/�~��=�h�>IT>�v�=�5�>���?�S>��>�yF>�̶�=��8�ID���ӾTdG>d��=mG�>�gԾ?��=]A�<+㌾Z�Ŀ����=-������\m���+����<׻�>��5?���6�>�:P>|@I?Y�e�H��>�㉾�p�>b�����ݽ?��>7C?OX�ښ�����l;h�=�L�>��?E�=� �w�<�C�>U��！�Z��=˸>��rM�]��>�E:?���"�V���;<�7>��>�҆����=%#�>���=�V���8�>�Q�>����>ͨ���=&H���u+={Ы<���>�s��#%�`J>�q7?Jq��4=9��=z�=�>���A�>5Ký)V)��c>�2y=����i7���<1H�>�ɚ�/9����ݽ(��>����$E��j���u������9��k�վ���J�=<�#�� �u�.>�!�_�>��ƾD��h]��#>�U?���=��%�=�yݾ{{�;I�+<��>Y��	�Ͻ�Zһk�?�$Ž5�r�>łh>�K�"����6>�e�>�m�>J�<��"
> [�>$2�>z��0�>(�Z>T�V>�l�o]��Q���RI���w>w���g�'�o��>����  �m�
���.>������O�û�G�>
c�$Ӿ��<�[>q����'>3`=�Q),����<���=Lz���Ⱦ~Љ����>Z����پ\���*��K�>��>��>k�f>#l���$���ɠ>br�X��I^�該?PZ������z��>���>I�/=����_U�Ȇ%>x?���~�D�T3�>�o<����VY>\��><�(�╋��|>��=?��?ڣ�e|�>v
���ᅾR)>>��>��>d��=r�>܁�>=Ff>PH\=�Խ�2̽���>h>�i���x9���->�g=��*>D΢��M.?�4���;�=���c|>�b!=y�����%ݞ>�Y���j��R�&��>�� =��E���5?�Ǝ��Ծ)���>���=�e����	�� ߾�� ��&����P>���>�	��7�پh�z��1�<ζ�>������}>��(=}J.>"�?�˺�	,�>�Ϻ>'��>d�
=�0�?y�=H]a>3��H_ؾ_��>}7�?����*���� �9��l�>Ҁf>``Ѿ��3����>�[�=?@�ݩ/;�_�>�U�仾��J<+��>}B��������������;fB�=�'?����Y<�oq��:?��V��c�=�'G>]��>�Ԇ��4>4�)>$�=)5�@�A=^�=S���D=(�>��?.Y�=��u=��F�3�#>W�^�\��%9<���v��;�=:�ѻm&��`M>AJ=� �����v�5>_s>X���%����<��=������k��=m��7�ʽE�u�h֘>��ڽ���=:�F�>�PJ�CZ<�D=b��>��ؽ)����"�����>��T=���=p��<�c�>�#��=�;�� �>5�(�1!0�Ǝ��0>�jֽT{�R	 ��.>e1нJ��<1ӌ=b���)ȸ=�'�>�<�>}w9�(>���=�!>O(j�X����W�=Ǥ���=%�����%�{��xB>S҃�f��9]�=�r�>}�>CV�� `����>�O�>�ʽ����O��>F >12���fv��C�>��6�zv���(B<w?�1>����񎥾�ɭ>���=�
���ýM�s>�(>y��>����Hd��X�<�;վ��d>�-'>N�8���о�>a�7<�Q���Of�H'�>��=�
��� X�$�=��=�'��� f>�?��E3��)[˽ϒ�>��*>u���Y���������wOk�+@�q�3=1�>(�x>ӽ-�ʴ���eL>>j\>�U";�I���=��z;��^��mp>�{��m���>�:l=--��b���o�9>���=��]�(����Y=4�=��,=�/ѽ^>*J=dF>�T>Q2�>�Ĕ��.�������/<Ḯ����0c��'-���e�7�l�����j>xO>��]��ؠ=�8�>T�L;,ip��Z���n3>45>�qk�jAQ���>[�M>m�z=�>f�r>��]=�/�|��`�Q�5ކ>u~>�>��꾦��>�i�=�t�=u`l����<\"Ž��轸G����ʾQ����<+�=8����;ij�=ozB�@��e2�=LK�>�9�>)���,D=M��>�,�>4�	>�.�A�&�beP��G�m�)��J��s�%>�v?�c1��?9A�^/�>x?Ƽ�n=����&�>{����7>�S!>����W�c>?�>�[F>Km����h>mm�=�#％
�C�6= �S̽�f���V=�&��?Q=�n�>�'���w߼�.�P7�>�p��uq�jź<�>�Y9=��.>h�S>!-�>�E�Y:�<jE��`聾ӵ�<S>G�>6�����=��=��<�'��Y�=��=���=�y��!��%���Ͻk�gM�=�!>~�><�l�˨.��r>L7q>kR��6>��cv�C�I���\�:?> ���iԑ����>�Q�$O��#��lM�>�j8@�!�V�3�S>$�`>g�!>�O�>n��>�ڪ���h�s�齯�_�O��_=���=��=h����kq>��K>�,�<�{+<R�m>ӣ�=�b�mٱ��`�;��>sB�>2��so>�l>=t���,	�.ܒ�or�>��=���m#s�J'0>��>����<�� '>�0ҽ�9^�${����^>��s:���A=QT�>�������>��>��I>3"Ļ�I�_����/=�O)=���>P�Q>��=�D��"��!�=�;T>.Y�=���}F
�My�<�W]�G֪=Gd�>p�<>�xK��֟:�F>��(���V�p��>���>؁O;�w9��6��n�1>W =��>y��Ѝ��(>�X!>��'�4t���u=4�>���	���ұ�;x/>,��=`'����=x,�=�;h>�l��������z>���=g�T>����R�>�E�<pf׺�j����]=�:��{:��b྾�s��CV�=��w=�p��ǽ+gb=n�>]�.� �=�}�=���=�����9�R�>�'�=��/�$M>� ���Z�>�2?e�ɾ��x��j��>6�>�0��z{�?y�-�>��:�a��=�~>�$�>z]5�5u����h�|O�K��p�?��wE>�<���>�>�; ��a�>/><"�����α<�mg=�=}V���`��Q�B�P=��G�>�jy��
:>��(񾼝� >DZ,>i���b/1>YqE���޽/�>���:a��>ٲ��N��=5�T>U�������a%�=�T"��F;q�/����>��|>����S�@�� > �Ͻ��\��(J���?S��@m������\a�>�g�=΄@��������u%p���Y���(��4I>��y>�g�>舊�Wo>d>�^D>��A���ؽ�$F��Qe�d!��$�8>��=`�W>s?�����z�����>T����ڽ��>�=��Y=��<ik�>��=>����s�f�8��<G">�����w��T>e6�=�2��퍾ُ�<���=0<�_9����=���=���->��=/P@�f�.�G��>Mu����E��C>IN��|d�%���z�]�RCq� 3�>��>��<OC�A{�=.�=��[=�bʾ�	?7�>G���3��(�[=����¾�㘾:[�)�彟�>�r�>�ϩ���o<p8T=l�<��4�ڈ�=���>�V�>�����<uL>�M�>}�%�K��� 1���Ͼ\0><*�><�>  �e�*>�)���DA>�J����K=�~o=���_bY���=�����<�>�>�}��mͽXf��&��>R���`O�Rh���Ł>8�2��J�B|/��v>��>�x�<'!��?>o��=�ꣾ�]ݾ��D<��=��������=�u>���=��&>�(�>vJ�� �1>��l�\.?��w=�WG�߳�Ŭ��`��lj?~=>��潶���о�E>΋�:D>��|>�L�<0��\�>k">|1:>�M
��>˹d>��,=�e����=`��%O��cG��n���Ͻ�E��.�>0ѕ���0>�Ul�q^N>Ҷ��f!>�ʁ>ђ�>�������νS�>�wb��V����y��Z=�5��=47\>���>
ɽo�*=]!�>��>=����<.����v���lW��r��26�<��>��>>�S��&�Q�C>��ʽ�B��Q�>��>AK�=�ّ��+��DZ>�2
��5=�U�Y=��<Vcj���	���=�T>�(V��xɽ8"�>wTB>��ؽ�������!z�<@�нՋ>z��=�Q��wf���4>l�"�'��>>��j>a������)<�J>+���mr�,�i�8Я���2���i=9ؙ��~p��顺�Gj���[����<�>�a
>��޼<
e<dm�=��>����>�����=���=�Ľ�W*�iW�� >�z��]��=�z7>�vi=9nY�d��ߣ<ޢ>�2N���žZ��:�>��>,w��<㘑>9N�=�.ξ
)%>��>f�>���G!#���
>#�<#&t>=	��n/�����Y>�΢=�6C�O=<	,>q�w�*�������]>��=�GC���'�J>��r=��0�;��<�	t>�(>�q�zO>s�&>�;��P��V�=����>�<�����۵���*���v���_�>��"��e�>���*�>�쵾���<J!�%�>��4�t��<?��= Nf>���>�ּF/��Go���+�>N��;���ҼDf�>��`�ᅫ����h3�>�>�A��ߴ= �=��>��>���>�Fj=����J2�H�>Cf/>j(�:鿓��q�Zf=#�<#~�]��<u��>��>�E1>��p��E!>����O��<,Y\<��7?�> �����о}�>}@k�$䠾}jf���>���=P+��ɡپ�j>f��=�K����Z1=?�Z��@����[8�>Z��<Ӹ�� ��!֗;��q��7����M
=�P�=��=46���=�t�=.S���7˽��>X"�>�˪���7���� ��䢐=�?cK]�~�=Z����>蟼��&=gI>��>M];��vi���5����=<�1>�x�>�c�A�N>o��>��A9�>��=wI>U�	��]���	<ab>�*ľ�ѓ�iG��b:>o&����$>�]�>� �<�U��/��>��>bǸ>���=�MO?��>%��>��V?���-��>H(�<@?���nV<>��Y>�1�>��@?�EF���)o�>,�=�Se>�����,-�����n��w�k>a�?^��>8?\�>λ�����>3߽ד?=����4�C��%z>��x<?#��>f���#����R>.:�=3�>2��=�@-=8^��\�>��Q?������M=�cV���>�PH�����T޾s��>	��>PH�>���>��R?�q)?�U,>łK?�H>��=*�Z��t�?%;d���c���k�=��#����>��a�J��aM;>*@�>�/[>�6�=���q��>~�7>y�ѽ�@���1�|�Ì�Iҝ�Ͷ��O[����4�I�[����&�=L&���~>X�,>����z���lM?��+���>N�оS߷=4?�ߢ�=#[�~�>v0Ҿu���Ľ�(?B�1���l�������>�1?����>De��q�>����C|�G���Q��
'>�0<��j)�&�%��3�>Y=���	��Z��",���0r�2��0�
�C�ϽV[����=��G�=x��'�>0o�.�?6�ɇ+�xͽқ$?|k��L:���fپ{�>��>�����Ҿ�E�=^K�>Π��,�>�����?�&>Bj��؀������^��a2�5\�>=�>��ռf�?��>P���C�>��+��">?���BҺ�|G>(��=�%�s�k=���<ͩ�>�&�=���>ݕh?c��>i,�<w�X=r��K��C��Y�+�XG?4R{��f�5�>[!�;�R�!�$��ZH��P(?Y l�lо���=O�;��?)/��k��Mf>��i>���>X>���>Ψ>ў�>�$O�,k���=�?���I>=�;/��>UT��W[�>��0~'=dtJ��屾poܾ���o>�K�>���>��y�f�K=�^>�{?Nw���IĽm]K?��>��	�S}>��M�?�x�>��>n5��V��������>%g
���?_�,��᤾�$�>�-�����Al��o�n^>䆽˟;�Q?G,�~���g
??yž�����%>��C>ͧ�>�D}��	�=�ZO=*�j����+<������<!�^?KG���Ӿ|wj>�o��U���7��D���> �~�sܭ=x�c> ��=�i�Al=W��7Ҽ�����7��L�M>�.��^��>�qa>ۆ��}�s�b�k>gv\>�=[�����;O׽ X,��I��d><��>ɏ��Y>�
��t��>F)%>�Q��J�������;�����P8=lKϽ��O>���;�rȽh}������>-u�>����=�Fo>�9�>K�>~��=��?�`D���.�`����˾ ǟ�;�K�Y�?�?o�j>��B={?є�m>�".?x�%>���>����K[=6�>�E=t��%��>���0XM?y+�����C?A�O>��Y�H>���
m"?��>e�=䇼0}@�
�~(>+����`*?vQ�=5�k��&??D����7?kuH?<�׽6�?n�)?l�4=(�>���3�>��u?C]����,?��O�@	>>:�>�1~��5ξ�E(��E�~q�S����^���Q��Cb�Cp3�2�?� ���v!?����)�?F?����e!���N=z�2=)ϛ>_��>�H>��)>)��<g`�>M� ��/�=(����t�>H����ٽ��>??�>)�=�mѻf�=ވ��s�	?��Ͼ�q.��?�M��>�>����P�=�R?n���g	b��r4=d��G���A�����J�fľ��޾����!P���<��>�6>��>�r>��
�һ�>���>-��=1��=�@#?q57=��>?d��<=����@Y�[���+l=NJ����4��JG>�*�>��Ҿ�4>}�,��x�>�kӾ��V���E���n���46��*>�8K�#;�=�՘>�0>��t��b?�=&pu=���rPp�?���*��R�%����=, *�-HK�*a>/q�>1K>n���x�>�+>�X>]`�=v���e��� �x�>?u?��N�%d>�ﯾI�(>��<>��C�6Z�>����9
���>O��� >z6��|����S����>2!8�K��=#Q���>F�>L�%�iA�=d?B�ɽ?��+�=jҽ.=����k�G�D��>���<�3o�eǞ>T�L�X콞����)�㍵��҈�?|D���m����>� �>�\?@L�>7�5>�7Ȼ�)���kO?�>��ھ&E�>i~^>Nw�>�d#�+:?�ʸ>�?�����>%D?��=���>jǝ�p|�>A'�2ܾZ��=*b_>�`��̆���<�q?*?j��>���>��>��
>W��>�N��|�>�55� @-���8>�݋>�I�_*0�K�-�>�W�J�>�0?->�=vv"�?��<��=Z�;�ŀ��mD>�.����=}c��(�`S�=���-9 ���H��TD>^1�`�=���N�>J >�x?�mt�ǯU=� A?9B�>!8�,m+>W:-�u�:?�`>�+>�s��4���Z��-�=��f>VS�>-�h��4��S�>Vi��6!�
� �u���@��>_��>0��>��3?p�=�=I�&=���>��=��߾bW�=DY�����-x">��>tT?�`b>�h���=B�m>G�>��O=¯� {'=�>���=��{��w��su�=ܾ��,G>�T�>�D�	�R��)
?W�?AKm=��6��>�r|����>���>�&�@B?Q�9=���>;(�>���>Q{>��>��>�mW��$?e��>t��#>�S�<L?�
�l��w'�uB��=���B���DF�t�7>��D=պq>U�d>�Ž�6?o�P?8QX��B�>��=F�&?���A�g����e�	?��}��(�>�9����>o�==�3>��i?][ ���ƾ��	?W]���>�G��4)��x=��0��-Ǿrʽi���30��ϗ����>��=��>I���L2?$��>�l=a���>�1�=�wO>��G��"���>�>%Xc�<��Z�><���)=�����>y�R>���5���ʱ���?��&g�>�H�=9��=!Hx>� ?ZQ�����=�L1���>���/'��6�K�>��n�b�����D����!��/�Ĺ;��4&��K=�����>j�}1.>�;?;km�])}>G�	=X�S����<!��%��Z�]�`ό��X{�O�G>�᏾N�ҽ{l{>5��>(�>q�㾨�[���3>��q>�oa���ʾ�x`>W[q��>CQL���>�[�?�>���]=@?�?.���3J�9��=��>=a�>��=ez�=�{�=�4�>�>���5���D�(`�>��3�f�Ѿ����>�>%����^����%��>&��<]&��'�*> �>�s��`-�>�)@��@�>�u޽[m`�P9�=��?��I�����*�$����=EBN=~�?-��������>�-�j�ʼ�[��?��*�F?�R��zC�>8��=g?��S>E2���w>W����$�>L�����sO��3�>��f�w,e�I�3���>Yy>Z��<�3=e�>���>�u�>��3?Fp?�1=)P�>e4O�#�>u�g>�9�^�T?���>m>	�)>ճ ���9=��?�P�>����5�?���)ƚ=U�þL/�>Œ�>����Q4�|[I?�G=���=l 3��ޗ>��s�0�4+�5k�><���k��8�
�u�?>D���=�)�N儾�'?	]���ޯl�8�t�������(���߾U?)=�!i<���:��>᛾.�N>ـ9��?����WT=oT>��Ľ�#�>A�M>7�'?� 2>a{��M�>pf����j���7����?�Ҡ���>Ծ�K>���>-�g�Ծ����S�|j >aQ��j��=2�=�]?ÒB�]	�=���Ng(��fn����u��ek�>�GM��g��ϒ>b��?���=�\�=�p�=q�?�� =�h�>%5?^�{?n��>e�>e�>D5��Mg>�z=��a�=�:�>"� ><Z���%�W�?��	?Я='�<�*�/�ܞ ��>����.?����|���S[����>�:����j]�>|q?�ː=�Z<������B�D9���־�6�=���|��*º�-��>���
>��>;b>�91�h��>��>�T
?f^�
$������B�=c?��ݽ7R>�{�>���>:2���1	��XD?���>E����V>,i�>�e3�o#����?�܎�1x�	� �XT��cҾu
?���>�T�>eݾ��L>N3�>�&"<8�;�\iQ��O��3�@�77��!.�x絾�H�.�>π����>�\W=�Kj>!�]��g>��ƾ#?�����׎�>�Yg����%=ۋ���=&I�-^�=Gē=��>#b��Ę�+ܘ�Rt3?,��vl��c&�OR��T>6o��,�;��N)�>;�>"S�Wǆ�-)�>���=ժU�Al����Խ�&*����-�>�l�\����,��ͽ�y\��l�=�q��lz>�����j��gؙ᷾?V�c�����S���q[��K!�~�a��j8�5?�*>Y�0>��ܾ�㙾�h�>�D�>Q�h?�3��s�d��g��w?�q��h�R�V���>_`��v�}�ٓ??y�5?󐀾|���`>���>�즾Ń��]�>pБ?�{�>F��7�z>#�U>�"=Z��?��.�I�w�2T ������3���_��9GM���?)�B>c�=�1�<�ۅ>رֽ��k�2tc��K?�?�>I)��1����M?q�?=��>0?�n�EL���=�`>̨>Vc>�[��,ϾαK?a&���H=������_��O��:5�q�Y��x��7T�=��>aL�>�D>M�>ߛ*�qٖ<�FN<x�>���>]$?����6�D>s,>�_�� F�����H�������{�/�>� �>ݍ��: ��1>�>���;�o?��R�=]rf�OϷ�O�]�=�Ն�g���!�#�#�=��>b��z B�'��=���]��<i�d�ü|�>1����>��A�q��=�Y�<o�<Z��m�ܾy�?�O,>zv?��Z <�纺&���B��:[R�	M?�Ͼ��#��
D���X��ԇ>�@A>G����=A��L >��c�"�I;��=���޼n�t�� Լ)�>��ɽ��?>�S�>Od>FY�"��;�>�A(>�ҥ>��=��ۑ=_�<eپQp���=]��<�[K>0�>f���^y���>�p�>kĝ�����[p>:�!?�P?�[�>��?��Z��V��֣�|�CF�>�[0�d�=�L۾����=^���_8=��>b?N�L=��>�C�����Һ�?٫�>�C?*���?X���ᚆ�d��;�>t��=*��>�Ӿ�?[*C>.�J>���^�>.:����;>\7u>��=@1�>�ᾕF>a$⽜� ;�m?��?kG�>?H'"���⾅˖�6CؾR�/?
'1>H�>ܔc>˟�K=?���=K+�>�p=?Ts3���ܾʰ���\��F���#?5��>���>C
����>�&=p�Ľ}0�Z��>�ν��3>Ӿ�?�Hv>:vG>t��>�ܾ<(8�6R��.?J�?���½ҽ�>R)?��	��;�B0>�/
?U汾B�:�>�Խ~�T=�9> ��������>��7>��B�;,�>J��>:Fپ}+�����у�-e)�A�>�iF2>��8���.�.e�>��λ�D%�x��gyH= X=�d��؆�> =?�/�>�� �]�&?X��>	+>n,?7�e=�|��I���E>$ɗ����f[�{�=��3�6"�=;'	?l?ۭf�LK�Ⱦ��׾�3%�'	{>��>jX(��9�f"U>��>Eo�����#���xO�u�i�8�<���>=��<!�_�'���+s�>J�=ȏC�+�־���=�L*��ᗾPx�>J�{>J,>�;;��4�>�u��OO�v�D�ڽ�=�Z����I��?u��=Kt�>���<;���]���.�sӾtZ>��v?i����A�tC۾�x�<�{<o궽4�=M�=���=�l9��.��<?���q��ğ_=�1����<ʐ����ۑ�>��r=� ��V��	��>ͤ-��W�>s��^k��M��:%Z�e�Z����?�8�>�M�>j9?�j ?�Y����=��>)�<Tt���ɾ��I?��>���>!��>f�	?l��>ʜ"�x�ĽP&��?��&<s�#k�>��_?�_��7�A�حE>!�=,%���}[�=ѱּ�A_>�q��R�?�' ���6>`S�=��W� S��]�>z;��赚����C¾�o�vQ���Uw=}�d>�=�T����C�	A�>��>��ʠ�>�E�>�>��׽yH��j������i���00?�ˎ>8M�>>׽�d>�������=Zm��hl�>>���>hV�*?~��>j��>,����|�P_��:�>4���>�w�ǭ��>=�>:rN����>���>�P��A3��=!���*�;?vˑ>̢��#?��>�֡�c<���9�>�v�>Y��򊩾��?Ђ�>�<�>����?|�.?��Y�>�=2�<3��>[���Q����>�E�>�X�����<�т���?��p?�O�=��Z?�<?$?cR�>�W���Y�>�?�����=Q��>�j�<��>��ɼ��м
��>;�*>���=�?���=�u�;Po`�3T��'���薾>��+������c��>�"�>���?���,�)��5оI,J�$��=�		�z�c=��>KY����3>����r��>7�U�ü�>a��>��?�E�k/&����u��>���g?>o��=�2O��Ež��5>Xl���s7>�	�=�˰>��e?����<��:;�]I�'*����=���B?�y�>��j>�bX�3ǟ>#w=�`���
O�S#?�����=������>-�>�T�>����:��0��蓾y�a��p(>�ۘ>�pn��ƣ�m��>�$=k��[Rľ2$��.�>�p ���?F4�+7��U>���?���5�ɦ=e�Q?�R�����ȝ|�'��>�'�ؚ�������b���0>q�z�Ӧ���*"h>E(�=8=.��)��F:��W��Wo�>��1>[��>U �>-�F�U��c>�oK��|u���<�!>�>�{x>c@��E|����=�_��W04��#<7 >5�*>�O�Qc<gWj?��>x�=:c��${3?O�u�p����=�
Wo��0�>x7�>�lþ:�N?	��>���=��?��@�� Ⱦ���L�(?�پ$)Q�Oc�=��#?2'��vͻu�5�
��>�7�$Pž�â���?��e��������I1~>����2P1����=�f5? �U��Gc����`�	>HI��:������>��9A��v�>�=&y�=c��T:*����>��>�)�����
s��˻��}�ty�=T�a?c��>�Ͳ��偾�+C�F� ? C�u�Ȼ`i�<��C?�ߗ��^.��#��%�?ᄥ��i����=��G?�Z�>rԄ>X}f>Y?X�>��>��>ڜ�=��<�I�=�ۀ���>I��=˝���'?,?�%<<Fb�>�y��n#=��n=�1;>\k��Z�����-��녾,���>k�� �n����?�;I� ��3o�� ��y���A�<~�A�/>�����C�ﾛ�C>-��ʿ������������cݾ	оC�޽,� �*�>�LO��"<�w@��w�=���>GRq>�H伦��=	7�E��>�?�"�>��#>��1>Ј�������>*S=�����=����H��B�=T�j<��j?�n�>��>�?qX�k���#�ٟ��)�
����>s�>���)ꭻ�r>}�{ڸ�Ym4�[�K��U?����O��<%3z?�y�?��?�P4>�#|?�(�,)?�����?��=��R?%>9���`��E���m~�k��m:H>4��>�]��W�b?a\�?!i?�w�=�ܾ�$�(��+���{?�z"�$I?�QH��F������X���$F>�9R>��>;~�����><��>�
��ۗ`=	��ay���W���P�:VL?��$�É>#N��I/>��A��@�=̉�=*�?�]
���=�kY���?�#�>J����=�?- �>}˾��w���p��%˽;�x�b�?aOG��J?�x�=Y1�=��<�> +>YG����޾��ھ�3���F>�.!?���>O|�>U�>��T?����'�G��� ��[Q�I�:��FA>F�M�o^ܾ���O�=
�?�<���%v�>]L��{��V7>��>�J$�G��>A 齭K?�#f=]���'�=�N?>��U���󅿷߸>��K��[���1>�R�?^�>6X�F������ �o>����5�!��>�է�+��>/�9��A���Ng�>�S���#Lɾ����g���;�>�J�>�~žG�ؿ��}>@ b:�Yi��JK:��G=F$]<c0��iĽ	{4?�L:��1g�B���\���>Iď������ᾖ��=�j?�&�> �>�n�?���>����ƍ���f���=�X;Y�1>1��@���%�))��i9��(s�_�?���=�>�`�� ?�R#?f�m�� ]��.�#�>n?�+ ?*��>kȑ��QӾ
*��(�9����>�>)��>�҈>�?by��p���5���x�>�ԾRdw>S]I?*W	> �ѽ��_��Q>�~�=P���iӾ��t?6�?P��>nD?6�?��5? %ǽ�;?�~�S��ͤ��ֲ��ӧ�?A9=R�%�~��nM��r<�7T�b����b=�羥S��=ฉ=�Q����~���?��>Z	�=�3?}G�=Bʣ=�����P��=}�+?B��RN�Q��i�Ѿ���`Cv�7��?��>Hʉ=X�~��p,=Gմ>����������X>�?�E>��@֬�>�����?���A2?F���F�>=J>��>����gc���4�WH��k�^\��x^����>�>�?x}�i��=����c�>�x\�a����0����D?��f>�6?��#?��?pl6��B?"��>D���B��>r�>d"?���>F���FK�]V�>0�A���۾~a�<L�l�;򉿽�žBa:>����������$��>�|?Z��@_�>�C>c�k>�����m�3Ҝ�1�žu��=�b>�Hr���=ds'?y��>{i�9��ŀ��������,������>g�^?i�?�?��T?Jg����Z���ꆾ��0?V��>�`�?֭<?��4�n��>����I������N�>D�5��PB>e/��3<���>��?�ȸ��Q]>��?�qi�	9��P�>�Q>���=$2�=M-?�l�>�i?�啾�����L���Ӱ����>�?��@�?���>�d���
��o�=-p_��/�>9E>0ʎ?��>��4?�2߾�I�>Q���(Ⱦ���>��%����>���>	�?3s�=������<)���a��>4漭?U�i?���?��n=�ٔ>n?�R���l�Xq��p'n>�����پ]��>�e�>�\�>K�=C���u%�����-�8>��� h��>�=z�l>�ҾZ?<?�3[�_�Խ�����mc>�x̽��پ�9���(?2��`V?��D�_"?F��>T�=f�C�V�#�:�dl��x4���}��8>��k������Y�>��/?�w?���>U���徳��>K#$�����U�=���=s�����ࠜ=>5`>�?�Z���'���'Կq�?���X��G|���i���>�6->W�ü��?ޗv����)�ߢ?���>�RU?�6�?�w_���>��l>�����=l"�=��6=�Pѽ'������>���˙��-h�>��>z��?�*9���K=CDξ0j>�v ��t=��x�=oQ�=�c=���>J��>+��v|?W��>A���T�p�x�����p�>�?�>=�>�.��ٖ�����ꃿ}�>��?�h�>��>��]?#�S>�nx��G���$>8)"���=Q�M��ą?v"�=��<ۡ��I>��̾t���p���婾�!>�!�>�C�����Q:�>�Z�R�@��5X�����Ѿ��4#�<�r�>d?�<��>�r��`�e�ZD�eִ��p/��Y>붉���?�?d�o>wkƽ*�?4ǔ>x�6��}><j�?�"��g����z�{��>,��=��P>��վ���>��?1=��I�lo��ߌǽ�3>��<>ȑA>Q,~�d��E��d@.>	�þ��>��?\��b=����>��i��F�?�%.=�Me������v�>�V�Ȟ=�:w�4@0?���>��=�O��� ��e��ؓ)��>���Ѿ<�����=�@B�n��=�6{?�Ő=�f
��>Lݩ>���<O��-?)�u>�-�>�,�>P�J����ax>����,�=~,��Aɾ�MF�!�>�D6>�M�T9���jK��{f>�Ƚ�1��s��g��?���-�]��J���|��X��z>��W�|X?��?j��A<>�:H?���>��|�v��>X��>q`��	g�=p%�k����ț�d�ྦྷ��¹�<~?A��>&p?;*??��/>���?�z?}x?ä�>,���EF�sl����N�?����07)?�	@>^�>b��Ner�<�?���ϖ ������/?����˚�,Tb�󁕼3�>ln>C�c�kHȾt@�a�z���о���^d���W��>?�Ы��'�>>��=�Z>�.���{>~�����>P��S�>#fh=#u_?�#�>� ��y:?N����>��.?��>)'�&��>>��>��s?�]a>Z/���Ii��=�[a=��L%��(?�N?��?s�= /?�^]?EΙ����L�����>H�g�=���s�>��?F��>���u&�?�l�>�/�ܱ۽�%��D?U�>G�d���T�>#�>�=P��l*�ˁ�������hB�Y͢>����S�& ���u����u!��kl�>�0>�e0>��۾�Ճ>�?�>��,�̾���������F���^�Q���\=O��5�?uuk>��=`���Yp��Ȥ�h0��n�=%�=2x? .��e�?&�?�>#�'?���=�L5?`ҋ�����x�8��s�>)� �Įo���>?*�>�M��w��ft�n?ڏ�=��e��(�>A�?ܖm?܊��>�?:;�=A�$�o�Q��������>�o��F�<7�ھ��a��x׿�' ����Gj���>�>i�a>:���C7>㸑>����I�������>�������翌�ƹ���S���R>���=�>ٯk�~M�=���>�����4Ǿ%�����??�#k���?�?3��I>r����;{Ѿ/����x��ۈ"?ݦ� ��=�b{>�x?l>�SȻ���[���#�>�w�
���>ZP�
�">N_ý�H��h�k>�e�>�t:�OT>M����c�>.??
?�1->�A&?UG�=2S�-�뾺�>r{�>�v�>3X?��6?t�>��B=-6��
>q��>1G������O? W�<)��8n�=�W_?���7����C0�|�|>�=��{Ѿ��!A�j�?�l���hɾ����=��D=����@��T>�.��������U<�-;? 
�������羋֗� Á�Sz�������r ?xcW?\�d?�?��?T=��Lg�k�'>�t;NhY>��a��{>�",�I}/�$�=���>]�w��(?����=���E�g>���K ������g>���g��<�z? N���n�=�\>�������y��W���0� =��s��7��IӁ���? !�{�U=k�<5�{>�ļ�\H=��u��`�>��>	�>o%?>z, ?��x?��>�	�>J: ?�¾�(�>;>�>�����)?�lf?��U>�����;>}���X�>Q�?wc%>�l�������81���7彍7~��k?:��eQ�=а�>xț�yM��77��y�o�=��.�g�q��<�V?�oC�c��>�_>έ�_rv>�έ���>��۾�U��Y�D�P��>�꨽2�軄�]t�Kڟ�ջ+=?�=��> n?:t�=��>o��>#+�ß>�[��=�q�=O	�=0����_�=}.j>��}? >r�>+��>�s��tM^?I��>n���Ƚ��M�#m ���=1[ ?u�> ��=��A�Ʃ1��;���?������>�M��&੾3��=�-�>�������<%�?�ݾ�&����>��>#�>��@>�A<>�H?�<�:+�Kn>=;o>O�t�R	�kx�����>��i������Ӽ�K?x�2>��r=8y�=Y���$�8��%�#���m�0�$>Q�5�od+���>1q_��� ?�������� ���̾��;S@|:�Y��̽�,����>�6<�{1���!��^/�m��	
��L��s�1?O��oᎼt�=f8���#?Ѱ��9k��U����=M�,>�I�=z� ?�,`>�u5>8�?������־��B�����x>fU�\h^>Q=S>��>�f��0����\�<��=	ƾ�wo����>:i?N���>�=��?T��>�	?{�Y?���>���Fy�򐹾❸���������>�Y>��>]d��ܤ= �=���>�:���H��]?��+>�����ԓ�~<>�ܯ���߾�柾�Q?���>%�?C�E>a4Q?��g?U�e>��y�Guz�X�;/��F��=�^���������*N��􆾤�3>N�>	� > �>��?�J��?���>�,���#���JU>�w�>AaD>�M�JU�?$sM=Dw��xk�ўW>�9�=|y��V�ɾ:*�==���j���Խg�֫=M��>r�����t>����؞=�,��q5>o�P>�i1>�&�i`+>�E�>KV�>��P�>CZ=	~���.&=ByN>ԉ>�'����U�Ua־C���N9�L|�=���Ѷ">�>B����b���>��>�>�X���	��(��p�>��?ә�>4�>k'�>�����g�>�->�����ǋ9?;�˻j���!�Xz�>bK�>襩��?���	���6���D�����U?<����Ț�L+����0>�[�>���<e��>w�>���=6Vi�c����CqA<x"��2`�>�]��j����>�>F>�~<�;�l�>�o3��Ig�p����,)?n��>`�@?^o>��>>��1�1��>�_�}����>�͠>��><��+�>�W2?��������>��T>TD�<+x���þ�a+?�Q�� 2�q����]w=1��>��>��K>�:.?��}>A��=�}�O7?��(��iսS��i;��"��k0��f?�o��f"�>!�v>��2=e��?�b>�H�>`e�=l����E���=�>�
?�ϕ>e���?�,�L���M>�w?>k�T>���q~��k]��+ k�y{=!E>�pl>Z��ˎK?m���k��=y� ���>v�K?�,ս����+
�>�ܺ=�#==�ݴ���&?�ӑ;rk��G>>�LF��8<�<o|>uþL��C�>��x=3�Q��6�S>�,�>�0þ��k��WU?b���#]>ƕ�y¾��#>�u=]p�=��꾚� ?�����>u��]���Z���R�y�N/�4Γ��a	�X᳾��>rf�>Jx>�iO����J?c>N=Z6�I 9���	>�!������1�>�쾾� E��b�>�jE��T%�:���Pn?Q����f���I�h?���8����.L���H�1�}����Q��^"�>�]����>Z߬�P$�>ׅݼ���lĖ�4�޼��>B.�z(�bm�!��I޾�#��D�_>�P�>��#=�'*��4t�!C ?o��=�$A��	��j`��!���]��Hv�5�T?1��?���>͐a��8�>��^��.�=\Z�>ќ��1Nپ��Q�і����>`s�=v�=����/���v�:��>	�y?W�@>~v��jSe��J?��d����)=��?�Aٽ�R"��D�>����+?����k���3z��zR��g�&>:&����V����V�־���i�O��罛���8߽*ӝ>����T>[ik>�  >�b�QA����>	 ��M����%��S?{�J>��9��.+>n�%?\��>�1��u�&�=ذ>a��8���B��I"h�����e!��b>��J?�菾�F>/�?PÉ>�8�?�Ny>�|f>@�;� !��%½��'>~귾���7̂=L�ɼ�ՠ-�d>��
>=�h�>3�H>�z���?��#�g�s��=���ã>)�4��V��<ɾ�Q.�Y{�ub��i�<�
��OO?]#>�>�ks�5O?6�V?�[>�v?���*?\Vv>H]���h{���e?%��>΅$��q=�i?��gM�>��ž�T��aH>]ȼGO�� ����Ҿ�綠���>�L�=x2?FH|>�F!�y��<�Y?PV>|F��2����=�u�T�����;"?,?���>�9M>�4?o��>'�.�r���
>���>�2"����=Y�H�4�h�о�o=O��>��h?L@h>+Y�>�7J?q�2>㝒�l�v?{�N?΍���?͋ھ��λ�E;>N\��F?i׽����>���=ew?`౾���=�r?z�=����黷�[����tp8��c$?G����M>��	��g���n������gT��y�?,�%�=��]��w%=�+�=��~>ă��C5=��=��ͽ�n�ٱ>>DN=r�D=$�>�{>�?�>;y7��о�U>Ո8�Į"�:��>��������9!�r����ξ3]Ƚ�����>ґ��jU�=A5$�j^?-�?e��l���&>E��=쏧<�����\(?zv=b��������p;? �~�uS��2,�kh�>|�>�sU�h�.<��>F'�>7��i�+��͂�w7��&;��U?h=���>�x6��3�>11�G����=e��>{R��9[���~=@�>�:�C5��ܩ>����Z�D�Q����<�>�7I�%�I>�l�=�o��[B2?���}=4�Q�3+%�9�ھ����.R���>����֚�R������>���>�����鏾�&�>�|�>Y��}�ܰ�=��=��O�E_��K߲���!=h!b>H��J�?$�>V�>ʡ�}�M?�N#?)�=� ���O��tž�@���r>�j4��y>gGսP��=I�ҾR�=��=��>�7���`%9�V�O>��0�NL=澤>�n�>t!�խ�>ו�<vg
��l��#	�����/�=='�Iv��2���>t�,��W�=�L�>i�Z?~I�z���3?ր�DO�b9>���=2:5��*<�s���?F�o?s+�>q��>��[>���>�O������V� �>控�u������=�T>~�z�q8y�3�>]�@>kyܽÀ3><�4?�M�>�;^���,?�j�>�4N�{��>�G�1^ڽ��=%����O>�&S=�b>����4L>�<�����>�F=C��=? ��x-?����(�Ff�T?�ez�G��>:a�͗��#���t��C�７2?�!B����{>؍S?-�Z��fj���>�a �50���Jt<�o�=?�]������>j� ��ھ�����V���<?���`��S>�8�>u�?;����0��yH<����=��=#�=�Sz>Na�=�6�H>޽(��
u�=���<��仕x�z?�>��>/�P=y�$����S�>�r���¿N���kQ�>��?����Q��v�=]8�>|�G�#���� ﾧI�>$�e�#����^���?̍z?�L�>�??i��>�q?�>6�?x.�?ǁ_>MFv?�J\?۝��^a?��?���?��/?~��?uV�?��?t'��L�{?�ؽ�ы�%%l?}&�=���?�ܔ�S��H�˿���quM�4j�x�E����q=����?o%��EؽjD�f�ӹ�mt׿$,n����>k��+v�?G�(��.:��O��~f�Nb#�����y����3��L?�D�@�>�����?|�>�i>��@?������=�*%?��	�2CP?)7I?@7?zj==(?�U�h�>��A�3�&?Q��ٜ��B�>�E0?#29���Z�	�K?����aU��0?a�+?�Pk�*� �@@�>�g�?�"���h������e�>��I\�%Կ�O0���s�A3?�F�>��ּۂ]�� ���`�?�h���i?�����c�?縰>9���#���پ�T���(��&��?RVz>��=�𕿼�?�wa>3��[a�QE����b?e2�1Э����C�B�� �)y��+[���E��셽=��@��9R���6?��x�-�S�e�I�����d��9�������7ʾJ���^���Ǿ����jj��a��\�6u徑Ž���~>���<x�����,P�?LU4>�J�?��@}��{c?��>��1?��<����h�u?�H��Pv�
g����o������ۜ�ZȬ����>{��>�὾��<>��|?y{?8�;�������?K?��Y?�� =z�>9W���?vE����?`iP?�#�>�\�����u9�M�ſ!H<�:>(��>X�쾉<3]#�}p@���	ֿ�6?Շ?���'y����>�v>���+1��}�?���?�Je? ���?&?{쾘y�壄>�"?��?��?z��>l�	>�����=���z��������>]�Y����� |Ƚ�>�.�A���a>����w��Ƨ㾮�#?͒E�H�tq�>�^��{u����,�*�>�v�>) �l߱���8�qo���_޿�\��T�>�"?��=n:�*�?Pp�>�DP?h�?"�k��a�>��?�А?2��?j�7��d?�{�?I�>(�U��Q>fD=ɶ�?c� �xa����?�:��^���>��oD#�	`�?}ɢ?K���%M2>��[?�2þ���>]���.�?4�X?(e,?U�a>�/ ?�X? �?e�l=!�;?7SF?GȪ>R�=c�~��@���_?$�?2����r�i��P[>�?��@3<�?-��?�ؤ��ܽ>�?�.ɾ�E>Jr���?���G���ӱ�ڞ񾦣��N�r����� C�!+��.�>˄|�2��W�W�n��� ���\�/Z?���?��z?&C� �?1A�?�eѿ�N�+�����
?5E�>yj? �>�.4�9Kk?�(J?�T�?���8�/?�z4?lR�?@ˇ>�~?|UӾ�N?�d'�u@3?�4?��?6z��@�>�?Q(?&Խ��T	?1�>��>�\+��Q�>m���BT��<�� #�>O�%���@��>�!@���?���>��/����?���?bE?6�?^����?�� =��׿�*���O)>Q9$?�BZ���Z��a��ڀ[?�<0>�F?��;=��T?�cӾ�Q����<��#�L�!>{�"??��J?���O��>4�h?�-�>*��?$��b�,?K�=6*�e����~���=��?�e��<������D�>Zu=h����M?S���S��?n��I9?��ľ�y�&�N>"t,� �B�L�¾rX7?�N	�V�>)}@"ã?��/����
�̾��b?�Q#���>�29�笠�M`��t��Y�'��>&r�G��>�*�?U��?
G>W)-=-i=?���=�=0���Ǿ��{<�+?��!?=��>R{	�������U?�,�>ܧ���ͽ��?�,��2�)��/Ͼ�aϾ��ھOɿ���W���N">#������f��?u���VVo?t�������X�?\o�ؓL�a:\��v}�ыӾ��������߀�h����B�O�>���=���?��;�B�w��>ڄ޾�ɾ���>6pm�������Ѿ~�?j3X�������b��7辛c���Z�"�I럿�9!�B�����?u�~?�?sq�=�1?�?7��=?n�h;?�!>�P�]	���>�O��|K�Z5>&풿�#r���a�4���ύ���!��S�?+��y���[Q?�W�?�����I���>� ,�2�ƾe�?M.~?��b����>:?�>.�>Bx�6�K?��<V��$�|�}�W΁<�a׾�X-�SZ?ݨᾲB�����B�=�ӽ=�q*>�>`7>x��,��`"��7�?r��>X\?��?�җ�W&���9�?oڎ?[	x?ݔ1��Ѐ>�#c91)����=ۂA��B����Ǿc�|�n�俈�i�� e���O?�0�>M�Q?�����q0?�rL=�?���秾)�+?�
������I���=���?��z?�`��E ��_ʵ>L.��=9�>�G�?�9����?	?��?�dq�{�=��?�
�ⰿ�R��a�%�{����y%�q�1���>R�%?j.��4�ɾs������?r�?��7��Y<���=�j]=v�ѽ0� ~ҽz��=IU��-�i��3�>[t�N^L��|p�u��>c��>A5��X���Vw?p�y8�%fϾX�M�j���	o>��?>�
�I~��GL?9s=4s@�@��l>�"�?��i?#�?���?(�?�n?l��?�LQ�G�0�=�\�>,a��+/�<�G��˃��I����N?k(I��X�>�
	�zg�>����"�~��J?���?;B����>�{�����pHh��"�<�k�>�j��<��ἢ?����62��No?�AP�{��>nG�>te�?�ڔ�Q��G�8�?�N?��L>˕<�U>�c>���Q�E?��q?�%">D�����(��F�<�V>lh��
@�;j���~��q�bܻ�`�Z>����Y��C��8��Դ��_Q?�L?d�?,m?о1�0>�\l?�\?O�?p�羾G�>�#�:�� �M�%���.���*���m��N�?�*?@��=�7��4a�>���?@��=~���:=�d?�#�H{����>��$>/w�<c���"vZ��Mk������Q��\��ąo�029?\��=6m�?HҪ�<M?����FJ���}���Q��?�=X�� 	�>���} >S�=�h?L�d=����rs�?�׿�g>Ey�@=�=ڇ �r�쾡:4?Kt�?XB��璾Zֳ=�j�?�5�?��o�"�>sD�>=e*>�t�M�>?q���/��-����W�\�?&o���4�0�>!/�>WLk?0j��裿T�U���h>A�>L$�>Q#�>[^-�0܃���}��2����P�}�9�x�m�hP,�r�̿>N?S�ξJ��>M�:?�i"?�>����L?Uo.�Y+>�zU����=0��<l�$�r����뾍�?��>�6X>�o����F���B>DA>���Q�ʾ�l?�1����=*�Ό��>)�쾻0����	��)н�5��;��-���%���>��>������K?X9��Vz�ۏ�>oG;?���?��6���>���?�W�?�U�>��K?�kd?)|>�d/�>Bc�/m ?���X�=h|q�p?�����r�>��R>>��?T�@`�?�l�>��=/��?e�/=��S��>
�w	��l��~�ۃ�TB�<�M��,���T��=�����%��س��E�x;ؿ�I->?f;>	'��������u�J�?�.
��Jh��Ǿ�λ������'O��VҿM�㾴IF����>vP?�O��^I?!�A�3ڰ���?��{? �9�Q�1?1Ы?ļj?��J?˕�=�d�pž�=o�;"ܿ��H?�������?�W�rW��St�?I�׼\R'>[�&>
�M��0�>���>K���.^>?��������E�<�����ξ���>&bԾ˷���j����?5r�q��A?��>C/>b�f=�!?�$�>��<rm_=�s�>�Z/?��
?�l>��>��Ͼ���=o��LR%=L�=dW�>i.�>00U��V6��L
?)2�>/G�>�:(�{K�gh��KȾ�'�>���>����?#�	?����V��>;h=��_<WY@���o��F�=�~>����FO��eW> p	���a=��=�΅>��Ⱥ�K�>�e�;ⓑ>bP���D׼�Ú>���>�ׅ��^J�(���e�>R�>f�>������.?��>I��m�>���>˚�{�&����=��A>��=w>����R?� �kY.�j��<[Y��R�>_|�>�"M>i鄾U	����?^�?���=��	��G�0Ƚ���=H��=�:�Gy����=AJ�j�վ�軾+�$>�l�оȍ�� �?nJ5?���f�U�>'��>!�>uՀ�����ܾ�W=�o�n�n_�>bf�����+x�3��<��>0z���Î��)_>��*�Q�>�K��ƣ���>�k�>�M+�c𣽁�>5ț�mK>�����g��=�g:� >�F
���Ǿ23r��D >d5,�AR�9e�r��(���%�̗A��V�p�>[0��k��2/S��`> 7�C2>��v㾒�? 	
>P�;�j�=>��>!z�<@�4�-V|�	���'�����>L=�>��[�,V!?Ҫ�>mMb�P��<���>��C>lA�>�����=>v�>>$�>g�T��@�>V7?.y�>E��=� ?��j�cMľ�t>D_�.��p�:=�(��>�i�xJJ�|%U����>Ύ�>�u�>�x>�Wh>M��=y��}]���-?�^N>���y�5�6|#=_l>
?�>Vr��h�>G�E�� ?�2/����.�?���<���[>��>-?��5������/��>�s�P���}�b�о�镽�
����4>�hھ>��>�.�>+>�>���=��3�b;�>�U>\e��$�"���>�n�8X����8����>b��Z1��,��>��򾛨�>S �>H�߾pP�=��>�+���;��4��A޾�X�=�!���Ҭ>ƽܾs">����=�&$>-׾w�>�X�>��3��[��f�>WU�<3~!?�=��ͿF���D>��?@?h)>���I���:��=tJҾ�����P���Z~<�Io>�(��Ɖ?�$���$˾�
���4���M.�o���M�!=K*���j>�t�>�b{�,�׾���=v"�<z��>�z̾݅�=����=g�!�i;��i�>z�> G���`�=R�&>�>���ݩ����f�?.:�E�z>���>��
>��>VA�=@���"�Ǿ���>�>��׾cB澫��Oر>�^�>k�>�%�>o����9�}���;���`Q9�\[�[%C��ߘ>g%>�<f�˻3>��<�Տ>In?�q�>~�	���{��x�<v{�>��<^��C?��+�>��;f��<m\|>s�>�P�B�
���>�;v>��2�D���N>�6���7����>j	P��?i�>߸#��'�>�\>���>�=�>�.x>^h>�u�>GΗ�oU?�
�<���
�"?L`>�E�>��>��о�ϩ>��(>��¾�q�
��l.�0n���.����>eG��J߽�,L>̕�K��=�?�H_�>d" ?d>$ξ!Ȇ>��(?_Nt=��?+p>��-�J�>�">=�Q����=K�o>��.>��Ѿٔ��_R�6Ū>d��;�C#���>;��⩽��N=����+� ?u��>ƴw>yw2����>XZ�>>�>�h���I��r���;��R������*���"�������n��=[��:����>��L>
�=����>_k>�N�>��H�ӒA?٥���"¾���>�}����>�X�dL<�����?����q�>1�!�֦���a=��=Wʾ��.�޽u�%�OK��k6����<IX��N��Be>>�ݽ�ē���
?���=�9��پMB¾�a���y$<E���櫾�ʇ>A��b@F���[>�,�=E�j�p��;Uʽ�Z����>�Nо�(H=J��>��)��=�<����{��躊��e����)��=6�mX�<���#>��>/8�;��>�Q�=�>��i��8�>�t�� �����o&@��i�>#����/���>ҷ�> �z�^�Q>��H��	o���?�| ���>��=��۽7�=�4�o�Ѿ>�1?zݾ%���3��l�+�����9?�7>���=*/�>��`�k>>�X�8��>��C>����!��>��>)����ԟ=��.�e�>��>@��>���P��>O�?���I�%>5�">�T.>��S�M眾X�Ľ9Z�>]ӽg�P�;��>�-�=��=����/�;L���?�α<����c}�����>=���ٞ�=t�ڀ ���"��'�[�m�O/=x4	>��|�&��>S�)?�Ƶ<�9=_��>N�!�F�w>Ow�������#2��'�����&ɾe�->�&�>WĢ=Nhe��߅><�<;]�>�;_��Y�<�Ȃ>��?�(I�K��>��[?&�>���7�=yS	>/8�0��>��>����$�>�9C�p� ��-�>�u�p^���׾��&������ ?�}>�u`����>���=�ќ��}+��Z�>��->2S��ĥ=���=_���}�>3�{��q�>�7�>�'>�ۼBj2>��>	�����>6T�>�p������u'F�%v�>�I�>l�нë?��?l�]>s��<��	?E]7�z+�}G�>����K4�>�F;=��>OѨ>|�>
�f��w?��>Y�Y��.����>��2���=�?�,� ���4����F>�I�=��E��ܾA',��������\p��_;>�a=��>oM=r$�>�6Q=k%�>,���s��=�m�>�ˣ>EH����(�Z.��G��>8����>R.�3��=���>.2@>j�?��P�*>�f�\?�H�>|@{>.������*���잫�B#׾��ӽwJ�>]Ȧ�hގ����= �(�-<Zi�s �>���>�=Q�֢�>-sN?H >��c�tZ��L�>�.��C�ܾD�O>�E�;��Ǿ2��ݥc>��>��𮽤J�=�8G��?)s�����>q�E>���9�>X�#>>�a���	>H[��ʟ�>��齎`���f�v�?�־H8��q���@Ͼ���:��_8��>����>L*��������m>��=8
�i?���>�#��I������K�R&B��#�=����������<���'�c���M>d�+=�1�F��GF�>�?�=�p�>�0�N���*�{�>�b�"w�=���=/q�>��,>H�'����>�?�n�>*<��ý�+�>q��=f�?��G=u鵾�Z�>`$>|�V��+>4����V>�E�1��1�s��>���C�.�I�>�c�=�k3����>�1>V�;�]>ڄf��S����<炚��ޕ�E�#?� ����w�����N�T��>���"?* K>d�ξ�w9�'B>SZ������e>��ļfh��y��9�5>� ?R�!?H��=J:=�n>�WU>�mx�g�����HJ?����)�gm���>s0�>fח�ѓ>�E�>��'?��>�G?��
?ڽ-� ?r	�=ڀ�>Pc>�>@W1��s�>n9���N�=#>8*�>D:>���=�!<>���>��ҽd�>v���W�A>�>=o�>�6\��?�.<�	$O��ܝ��:H�lt����P4��a�>�����ы=!���?p=�=-9x�o������>\~��7
��^	پ�b�����B�鼨�پ��\�o� ��໼I��=1��=�1����>��=M��>+H1>j�\>F�w�V�e>n� ?�����\=?��?{��	�^>4.�w�=�x۽���>�dདB(�;难��>�@�>���>�N?��C>9�,>���?��s�˽d�s�*����� ��4�U���`�>��>��?U_�I�7>�4?�Q>�F?r��>�i�=�e�>ip�>m�?�<���>l!�=m*?���>lZƼ����޺�?9:�?m?u+�>�l�>!i>�;C>�vE�z���?6��>�KP>�ޏ���O�s�"��ֽ�D>#�?F�����>#��?ˈ%�|�B>����_Q�������n\>e��>�T?�O�ӑ'���X>1���[o���=J;,u==�ک���>Y�P��t��!N?Á?[W,��	w�C��;Ri?E�>�
�?��5=!�"?3��?�֖�5�>,Y=z�[��E��fL���"\>����{u�=�G�>��=~��>��H?h͋>�н�g,ž��5?-R=�	����v>?�H�> �=�^
��þ���Ug���	�k-P���U��6����?h9�����`�Ⱦ���>��0�9L
�	=���? � >�7��+�=�by>�Y�S�r���"���?�Gվ����,M��3�>��ؾ�@��tgm���?���>���},S�)t?����N���|i�
9ſ9��>8qP�X@�;+�x�0>i���<&H�჎��X����`PQ�q��ah��z3@�������?务�P���	��n��}T���p���J�t�U?��W����'�x���Y? t'>/�?��G�G�J���+?�L��'!Ͻ�)#>���>^�r>�*ž�6���g ��:��־�8*>�S�=A5�\Jo>�_?[ń���=��=�%0>�`׾��=��=���=�WZ�+e>r};�?�dO?�l�>2�?&�??��2=L��>��R'n�#J�r���]�s2�T>����s>�ѽ��h�����t��=��+>����Z���ı>%Y>����#��y>>�M�=��_=�j?6�?¯?�����=ƾ1���w�?��޽ʵ��j(���6��=�!i>���*Y�>����)������r��G>JL�>D� >�O��K?���>�5w>GЈ<�� ?)�>C��>�?�[�4��/�">����ӂ��ە<v�R�����Wp�+��	�>0�q!Խ7-?��?"��=����R�Žb	�=R�?�<�>?�H?\þ��>��(?�><Z�O�Т>��A����W�߾D�=Ab�>�v*�81s����M{ʾѷ�d]@?�Q!��C��?k[?��F�ȗ��u�F�h�>O��D܂�0�?��>U�ʼ�?�e��X�6�r�7<-Ľ>���>^׾�`K��e?S����ڽ�#����?�ﳾ��?��t?T�=�q�>������o??y�����#$>xi�>�gþ��̾�$��뼾e���ǽ=����$����
���e=��j���X�W>*�=>0�?�]ԾM��b6W>��>��>yW6?ɮ>1� ��y���9B�� ��4�g<x�>f�����>{ܲ?�H�<8��;DL�>�+?�ي>�zt>pye�Q�h=	��>A��>��="��mӆ?��=$�w>�!�=(X(?T]�>A�>����\<D�?�Ţ>�6����8;>��0=�p�e�2��	н_��>rL�?�2>��>��= Y4?��G?zIJ�x�>䐕?dZĻ٭2?>EӾ�
��\?�����>���<��!�:Q?&v-?�Q=_��A�Ͼ�?�<H��;!��?~�j=� �7I�?Q���?37N�N?�N���=-���������^>Mk�>/�=���=��4��>�"�>�6p�I۔=֝��~�?F�c��[�<ׄ>��>r�=�V>��M��Y�>��?�,�=������;>����+�����`>'�Z?�E=�g�=M^���þm�w����F�6���1��[V��Z���#����!>�w�X|�=��<��?�>�B�<�F>,g�=2��<w1Q���?\�#�Z H���?)s<�wf�����vk>�7پd�(�9Q����>e=��8)�̌>|�>�K'��޾5�;3��m+\�,���=8>�#<G�"�T��>yQ��+�G?��>����I�˾���%�H�i=܇=�]�ؿ��>�Ә���Լ�.�=n�?��E>H�L�k��Y&Q��!�=�'��b?��>�&<��A�q	�>>�H>�ﰾ�Bn���4>4�#��}��B����sI��ɬ=t��A�?r�����Ͻ�+�?��?R����`��������=���h����>7��R�><��=�?�>J�7NO��?��.��f��Ͼ�;`���<�>4�^��V��tc>F�������uܾ��;��Q>&�6?n"�=�?�QE�>�B�=�h$�V�7��4�>�>m�����H��>�º����� �>�����>>ߙ����>Ey�?x$��X��<��ֽ8�B>!�����=3'>���>��>ӗ�-\��HX?�,@?�!�>$��>�^�Y��>�f�ѓ�=����wW>J� ?�?=c�!��$��C>�_�>c��>��t>]Y�>�K����>�2>�Ⱦ��5�����/ǆ>����>�l�=�G���󊿥��!8侖N=�~>;=�=)�}��Ҁ?:2y=��
?��⽩��>�>R+>���r�=hB<>���>`a��;#��4�������>��;!�ؾ�=�>�0��t
���>��=v��z9T�_�<jX?��S>��C�$�?��>��?bx���|����>)��>�/�fH�=߶�:��l>�ݓ����>
�j>�d��.�����"'u>MZ�?d�i��`Ž�(�=���>a��t�׾����o?��>�Q�?LF�=�m?~OJ?)?�>�;5?G?ۘd>e�� .>U�=!�N�z,�>S�E=�����A>$�>>��)?�W&�w9=X��.�|�t��=JO��������پ�v?���>	��������!�#n��?f���=1N�>���E�n>D~��0��>Xݙ>(�>ݷ龲�=�h�>�[?������x��Oy>���>��f�?2z��M^a>y�?���>���<Wt �]d&�ig?Q��>u��<x��`����í�`��<Ӡ�=:`�^��>1
&=�a��Dx�?�`��(�C?uK���?�3�i�/>�l��I<��8>�??)C�u(���?�)�[���>v?#��=�i�ݙ��r>�8>��>s{�e۠>K<t���V��5�>Ѯ�>�C-�_�<oab?�m���=�g�4߆��Wm�.��=Uӽ�e�>ڳQ�s��SE��� ��%�<�� ��������=���Վ%?�z>6��=�98?|��qQa>���<b��=#B#;�u����M��6?�]���Ǻ��O1?{F�>�丽| ���a?
�U=�
����=R��>;�=����Eb���j�?;@�>ĩl?޵Y�G�U>��>�}>���$��>�㨽�o�>�W�y�!`.��Ǩ���?�c�=��������G�>m����T
�K;��n	>�v0����=td+���>������P���>kɨ>CҾ�A��L�?Wӿ�L�;{i �G�"����N�ӽ��(?>rs�ID(�]���a��<ٟ��P��O4?ch>SL���t�>��>��M���𽴍�%�>���>\�ܾZ��>�0j>R��=H3}�9����ɾ�F�>�>C���w������H�>t�ža�������^�>iV>䨐>��:��.?hL�?��>���>�ُ?���<� &?:��NN>�Y�>Ó@���=r����c�?�h�6G.>�M?��o?��>~lY>\�>�/I���ǽ�0�ֈ�>z��>J'�7��*mZ>�te�����'���c�OF�}����<���?4ۻ�Dؽ���9*־l�t�SȎ�Жs��PD>܏���"<�X���wa��P뾑?�dd��64����rn�>�,�{�r?ּ��c'�>��c��`?�a?��׾1DǾ��?>��O?c<x>�ɏ>S �>�Ԡ�>�&?�Ǿ��Ѿ᤹>dh�/f>��c��<m��*��C%�>I�1>L+@�k�>�.>�嘾��ʾ�-�<L�:>�m�>�����<I��>����X���3�;@>�i>Uҋ�
�>�4�=��2>��~�W)?ޭ�=��>���=�9�>e�<�J>��>��]s@>)�=|��>���1�о?���g�>���=�>���>x'3?I��>�5�#懿��ᾂqԾL1>ǳ�>o��o?ם}=藹���"�O>���1�Y=��>!N�>v�}>�!�\ ����4<��=�f�>��>�ǿ>ں
�
{��긓=?ҋ>����~4�?�z��ܷ�1�N���~>��;bVq?,��X ?޻��6��=�&0�c�>d�̾ ��=���>r':?��:>>q�f�8>;��>v�	���>�x��\W���_m=5��>�W�)FM>Y��>\)?�%˼��.,���Ӿ�Y���o>���H�	��ӽ�h"?�n[�������K��?�>�BT>Ah������&q�>�k�?�X>���{��>��b��Y���.���9?8no=���2g�X4�=�"Y�;���-%�ی<?:"
?T�:��5�>$=������8�%�L�"=�Q ?|%�`I<M�нO��>��0�s�=걏��o,�;N>�#i>��y���8>�0�>C[�:w��k����=}7
>|_.��\z�N��>��彆ҩ���������5c<�3�>9w��#ھ�a�Jp:>�>�O�>>y~=j�!?���>�*W�=���H���8��v~=Fs>>�2��Ƿ�>y᭽8���$�*�=�a+=��ۼ�O>��>���>oS��L~���>�'>'3?��S���>^�><�sa���=bV?9�s=����K�<]=�>ØL?+Of>�;��-�_a>Ɇ8>������>
'�>�Qt<U_g��5+>$kԽ�/��r�J���<H� ?�%�>����{�>��<�H�#�sg�=�X�=&�]=K{Ծ|�ҽ��}�x�ӽ�w�>��=@���t�j�	�]0 ���>�^ �Mse>5�>u�=�%��=���=[B8>aIu��r�=�˲>>$?�ӄ�80�<��>�n<#=f��Vξ��>�!��a��n~A�O�<��r<���>���T�=��A>�pR����)�P���>H>D>�T����u>��Z��>���=��>����H�>�%�=�=�>��������>�~Ƚ��ľ%)>�<��aQ>7&待Ѽ�?,��[=��о�>���6��J ?��$>�\(��΂>��$?����N��4�?�����>׵E>o�o>$C#�,?ܾ��;>�N�>����v���.�ɼI�>����Ma�/D<���>Վ	��1����<��t>=-	>"�,>$9=�5�>�U��t
��e⼹��YK�[��=H->�e���l�>�S�>�~)=�U|��%>ռ���r��~�އ�=U� ?4?��7>w8�>b������̾�﫾� ��l��>��9��V���v�K�>m��=Xl<��j��e��_��=��<(S���zg>U̟>�l!��m�����=��>c>^<��������g=m�l>j�ܾ	�>�ʏ<�x?����h���]I�sK��`��>K��>U��<_�T>���=C}�p�����>��_�ʐ�>��=v
�=���<��J>��?��>\~����M�<z��?JS
?Z.=�d?C�)<F4E��ΰ�Bj�v-V>'eA�H`�=�#�>Mk����Y���)>�x?���=k��LJ����;�
����g�{��>���>Z�>b>�6�yQv�A��>�M8>S��C��W�;��<�^�=�=��u�=vɝ>1|þ�.ľ�|B=)_$>}H��0�>����cS�>K��0Ǥ>��z!�>�T�>���>C��~q��!A�����^޾M�E�<A�7'�=QM����^>��ѽ���>����v �=�й-T���99�u:�A��>a�6>˱�YK��4>?��$�(>�r
�=#j=�*l> V�>�l6�N�о^S��m�?m�w=���|����>� ڽ��G�4��ʁ����7?Tݽ���Ej׾�0�>���=�����'��������>CV�=H���>0=��S��>�#.��|)>lh�=1��>��߾��a>�_��8���@-��b�����>arL��8i�Hw��rz7>�Iv�~�F>��ľ�⚾�W?�8���k\�R�/� ��=����<?@�>#L<�2�=�u,?�5� ��B�-��1?R�<i�!� �R��_>0��-������K�u?��ba���o��t4��<��l�=��徘�ž���W���񣔾Dڥ>�?�7p>MC��Ɂ��Y�%P�k�R��!�>D>(?�X���-�>R?�����=4iϾ��e?&��������:8�><B�>�̕>~�۽y_>��E>qSW>�o9���>k�?�+���A*��>�_=Ě�="SA>ρ�>0�=;��_��gp�=ًO��TϽ�?��)Y����|�=������+׾��?Qf�>�:���\����g�����>|�J��p�>c��S�>������>����'��>�R�>�(>�px<7\��NM��������h�Z��;�>s�m>S� =LT���>�n�=�xj>�*澳 ��rT>d�>���\�:>R?J>42C?���4n���<�ñ��1�����Ѡ=>�N��3Z>4��>vԖ>���7����	���1"�>�u����>�����?�y�`�&=pI@�k�6?�h����ý0<��>���=�d>!">'�>�u����>@����}�>�f�lnֽ��a�>�v=��߾��6���ĽW?���>
�K?_�=?�>6�>��:fu�>r�W=�4�>�۔>��>���I�J���m#>��=?�=$@�>}�Ԓ�>^�I��ؽ>�hG�*з=�<���=)��A�>E�0>�7�>5' �	���F�����~�O*��"�@?%	?�X�>t �&/����>]�?x�彝Ө=��=#t?[Dx�5�!������8?Fe��/�R(�=����XJD�z�˽��>
�ȽM�G>k�>r� ?�
t>1e������Ƥ�*����JY�as�=%��>囹����d�c>}?Nb=]�f��F��pU�2�	�PG�s� ?�'�>�Է>mϟ�Xc��KH�>�D�v�����>��?�`ھ�e�=olC<�9�>�㠾�_��o�>�b>fMF�[�W>�	�=�{H��>�� >��?�q��{=>eH�=�׭�$Jc>q��>�}澱�޾~n޾������7�pg>Xv�����9=��>\��W��>=�����V�Ͼ�9��Y�>� =��zT�~Q��mԺ��G>$�񾒆�>5�@=�_�>.^"�?��+p�t�=X=������?��?�$*�9���^d=��>� F=�b�!��6>��>�茶o=�!�=���>Er�����T)&>�۟�w�;>K�:�D%þB��>�%>E]��hC���a��w�=��>��<18�='_�>���b��$��|c>�o=af
�b$�>� 
>�N^���a/.=`B?>�$v>�ﴽ���<��>j����5��|��oNc��?І,�d�>a���\9����¾�k��a9��d�;~��]%?M*��"�	�c3�>���>k�`>�G��@N��U�C>k��>��Ľ	�ﾬ<(�'>�'u�0����*��W�>�;M>dap�v1R�U G?`ݫ>�Fw�"��>J3�=�O���^> =?Bf�='�>m�G>���>`?��>K�>"^Ӿ�3?��+>cͽA=�o�>4|��J{>j�߽��>;�|>�o`���&�F?�r�k���Fዿ�<�>�e��|��{=��s>�wF�1M�|�t�euC>?�>�/�����}�>څ��-�r�:�Fݽ�;�TK��x�0��j�>�>��>���Q�h��>nH?����\*�uYý��?V��=�C���B�<��&?���"��>�[�AIA;̧
>>Z׻;8%�Әj>d��?5c+>C-2��`�>)�u>t��>�︼yޢ����=٢?2w��Kc�q5=C���o����D��1f#�Ar�>7#�Ҟ������\�>
��=b���!?eH>;~�>]��>�Z�>/cH?���=�ٻyv�>@#e?��D?>��>��>�\?W
\=V�j=��>ΧH��+�>	?���>�qX��|�>[��=j�%� �۾,�>�.㊾����u��>��>NIr����>Q�X?����6���?QM�`�>����gӾ<�=��.˾\s˽e/@<��>�p
?��_>�A��
r�>�:�'r>t���Ez����^<O�?�j�e����f�\�8
�>�k+?���=_�>��i?Y�����<UM�?^2��7�>6���X��=�擾u�־�q�=�g"?�g��0�.>W�%=���sW=]��>[�/?�þPo��I�>���>'�>����6���v��*���X��Ǫ��8׽��� �>�V��.'��)��PY�<C��HTl>�JA��ԙ?�&�>�v&>�����>��N���������g�>�3��ۏ�)K�?~��U���������b\I?�o>�����d��ܓ����6n�=[��i�4��\�>8?s��"ƫ=.�SI����>U�b��>�����Ѱ��m��q�=a���pX�>E��Y}q��E	��	9=�㴾v�B�Nbb�0?��0�K�lbH��e�Z e�a�>Lh>8�� �1?I��>�:�������0\��0�?1ϼ�Ҝ<�;�j�x�A�>O�3=.<�����>9��>U��4Ō�%z�>�����ؼ��o�.�>|��<����Ǿ�>�?���>�>��O?��<��⽭.D>K�6? g(�I>�gG�M�eNj=v02�2�;;��=��>0h>^�y>��0?O>?�i�w��<�?rJ�;A���G�>סi>��Y>>6ҽlN���>E� �J?�Dv�B���L�>g�?��id��ּ>�������>^�+>��+�����&*��>��]8�����#=��F>�>x�F�.%?��1?�u¼VU<k�;d��=^z{?x�{�I���#I�<���>&�������#�=e��=�d��h�> vw��u�n����������z�<?�C۾Ϡ�;G������뛐>½K䨽���jɖ�ק�>K�>U�#�D]0?]Φ>*=A��P��>V_>@�>8������lc?>����t{9>�R�=)��t���-?n���j��ѳ�����<#�Ծiv��o�sn?}�ؽ���6����W���l��=״�>_�򾖔*�D�>'���?�_��(�p>��>N$~��ľ����o7>1�ƾ�|�(�"?)��>Q�&���>�N����>�f�;�>�r�=��6>pG���>A0,<������?>�;;���3��m>��=�ø�&o�>�n�>8+�>�q>��<>[+�>�06��T�o��4�$��� ����)��4!��H ?ռV��{�=�K?���=�7�?\�>��>�uɽT��=���>|���8��,�\?��W<W���h����6<P�<?���?%���Ӽ1��>�?����}E��!���f�=�B�����>���=��Ͻ���>_P<.F�=H�>�$1?x.?�G\?9[(>�)[?��>~�>,/�>O����=�L?#t,�{@>j+�o����C�>3⾯l�9r�7�'�)S/�Ҙ�=�r>?����]U�6?��������4�p��k>k�?}}p>�ܾ�́�Q.4>A�">��>,f<R�;���>���>���2珽緑>vrV>�þ������>If>�=W��.�==J,�i�`���p>7�ھz�?j��>wP'?��7�_�?(�>i�v>�d���<�/u>9!��`�F��v�6�x�ʽ8���
���=��|�t6D���>>��P�=��Ծ���>���>*��>���?�
���I�U�?<r��>�@>� �<��>i��ɽ�=��R">��&��g���
�l�>?J����y�,�B�ʲ��[�&�'�h�r��AX�3g½ �ν�F�>�⬾9F?��>m�`=���1�Ӿ�P��9��i��FJ�R�?�\=4�L����>S����F>��>0>t�>��������{H�<�U�=�?=�i=H߽��A��n���C��0��8�þF�m:�0���AB�����a?.�>~�������"��-?�_���Y��2��:*�h>��>Cѿ;��M�BP?;��>�%�=�L)>mGY�!�>u??�V���0�>��:��[��თ��֐����==��=r��������������-?��>��h>h�?��nh
>�x�L?�=��S������[?�������F;�jÊ>%��>��o>�J8���1>ǝ??,���η��??�!�{Y;>��ʾ������Şk�������>�>E�C>9X���=�\ٽ=�?>� �=d@?[�]���=s���ݝ?âa��]"��<�� �j��m?>%��< ��>�ɻ��9�>5�M=0�?�ů�%�>�>d�N��k���F־	���|�n�ؾiF��1(=QxU?�'�j���e?j��=�'=�.����=c�<?��Q?*$q���2�p�Q?@'j?����}��>>k>�<�kΡ>��.�#E ��9�>���/->���>��P�"s	��N޾Ā+��N�>��n>�/V>o�B>��
?��2>������>�>�I3=n*w��2�<���>/�=?t������>̀��(>핦����|??���m04��~>��=��H=�<y>g-ؾ���>٧B>A+>9io>��>��=l�>d4?�f�
� ?p��>�x,>ټ>zʩ�O�1����<�l�<#�>h6?���>א�=nf���)?��|���?�=F>��->> ��^k>�X,�q�_>��=Ą�����Q~�l�#���ｿp�>��?,�>�l���!�>����	>�/a�?dǾ�Y> Џ?�!����e�k(�V��>ֻ�=��=�D0>�𝾮VZ?C������="�~>媬�?$�>�r5?H���� ��	��T־�n\�c�M��4�=��G?O�������?rcd��?�����J�e>�"�?�ӵ=85���Xs;�&�>=W�>��=��R�D��%*:�^7Ͼ�ݎ>Rd?<H�s >3+>�ϗ��ب��~1��Х>�?I���rm?���ό�2̘>֥�=�+D�	g��>�H����q��A���^�>%w��K�龕�a��a����=�B5A��N�&�R>"L���T�X��>m��F�=�?14���M?[������f����P	������κ��4�=O~�<��g>��5K�>oVB>��e>=�M�~�=�?Õ)?G7.�vs<����>�p�=�ͳ=�5��i>4��?��K>�r��
�>d�w=d1�>�#�^�mRc�(�H>scN?�G6��tH�AJ�>ݓ��e�
��/=T�<�/> X���Γ����[��>�(T=�����(�o�?�</>��L�qE/>�U>��w��ȼ��=W㱽�'=��D#�<�Z��5?��w���l>뾚���Y�>���E�2����<q���Xþ��?mk��(# >��2��:�����S���<��P?�?5h��,���~�F>y�=�w�����|��k?�Wﾉ�3��Q����>p�G>ͩ��b=Y?��>h�=>'?T>12<��>��L?������>mQ�=����?H�>	{��g��j,=#��>�dX�:Em�s >�?
Ⱦ�b�>�c����>D\�<&����&��f?Œ�=����78^��uý�������*L�G)1?��X��#�ub�=�'���N����B���t��o ?#C�=�@�½k��}��+����|a=d����M�՟���i��ڇ>5xt� D�=�к��)�?��?�I>Z��\%��?���A�>�f�>���=�/ջf�>B�p=�<�w��>��>P?�q�k���4��T>��a>t�>�d�6F⼺���'G2?e���qV�]�Ծ�}�Լ��i��RĜ>�;>�T �Uy�+OR�D	����d?��E> �>��a>�K��^�^>�Y?פ/>i��>Q��=��=�G�>�	>�w<�B��?6Q?��}>����'%>V-�>�y>Ӄ?�n
�=��=M�>��9?�x˾��_�9���WȾ���|�	��eB>;��>�?�R�=���;����׾#�w���m��>���d���.>���>[c�������ٴ�Dk�HPݾ�̢=��-?_�&>�پ�vd>�:?)�1?m���:<�F�&�]*?޼ >c�)=jY�=r�&?��>��ºG�f�B�žM-e��S徘 �=���> ���z�(��>U�@?��i=L1?�>x�H�'�^���t>Cc>��D�i�)>���>J�e?m?457��-C����������>M\��Uh�������	p>mM	>K<�C�R�x�O?�d˾q=b�����>��׻�~Z�,	�٠B?�"-�������[� ?�u���HI���
���?�4�H�r�A:����?�|>��\>J�.>�E�>�� ��p�a�?�Q����@?����]�>c�(�>0���g�>8�Z��&�D��-L=�1��	���v���?i�9�/�	7e��������}��� K����>gK�>�ש=�Z8����=r��>{0��41�l4�>>��>:�>9�ະ��z����4?��=��I��v*!������=����#�=$Xs>	>�cG��1׾:7��<>o�	���1�>�>+��>��H�v�1�R�=߲�>���>�^�=C��>�E��F�����Z�*��%y��38�$���?R�������>�� >�p�>�{�i)=��M?�k|��ۉ�q����
>B�=tVD���
�Ă���8�=�|Y>���>�b?@f+�U��=e��>,�h�Uq?d��=����)�W��wԽ�׸��a��|�?%k�<"��z8R>3��֣>I����$>�7��d�=O��>��>S꾀�G?/�?��R=☨�Jh�=4�=ȠI�V�i�hqt�O^��:
�/��4U>�%�>��C?�����=���>�
�>o��G�>|���Ż�=�>��9?�E>7_���2
?!��<D)��I�D�l�����M���q��8��b�=��=5�]>�?�O���*2����<� �>\9B�lrC>��"�������<���x�ؽp#>̆ս�.�g�=J�?�޼�v'?u,������˽C.�=�@�<}���^>-#�=K�̽�ꄾ�,�=�E�=e�<�k����>N?��s���w�NC���^>�� ?�gW>U��=�R�>6��>e�f�!��
��,������=]0R���@���*?l�B����:[潉��>�;�X=�H[�<2����$>t-�>F�>�?Ϭ���f��,�.�O=#!�4Y�>hP�>�X�>2��>t��>$ى=\I(�1�?fy=]�,�@0�oC9����>n��=�!x>>
w�㰛>(s5?ȶ^>�.��o?Py�?�퓽�o�\Ο���'��I>Cc��s	�=<�B?�b]��ƪ=��G��զ����?�P@���Y?�)�>�K���&�<��:?PJ���%����%���8?�Ҧ>f^I���>vm������*<�=��ҽP%�>W�?P>?-z���<C>���<��<(�{��\N�A�=Թ�>���8<�>ृ?V�E>L����<&?ϐ�>7���I��'l��h��>�y�>��=�:̾�I�=4P����>x� 6!�GC�=�3��f�;��m9n>:`�>E�0>�?8���̾��>��?'�A��>��q�>s}=@��>B�=bE�>��L>�B?�I�=쫆>��x� ��ʾM��0ƽ�YѼX䅾H|ξ���>��>[?�Y�=��/?��/�)�����=�Xa>��r��!��;�>d��X
>���>`t <@c�?Ͼ$�&?�<2����ǉ>,� >L�྆��>��>Wh&>���캥���>U�'�* V>��>�g?�Ȝ�ٛ�>U�$>���8%M�?l�>��?�$@��+���D��=d��Z(�����.�5E =S'�>?*��>�ɷ>Դ1<�˾k	m>g�>B���H}����?hs�s\��?L�?4�+����+?t���)D�>BY;���k�M��ܓ��
��f�\�c5�>6�?��о�b>��1���>z�>~R����?k��A�þ�� ��� ?,{��+Z�!��>�r)�`��r��*?�m�9>r�P>/7\<∏�;(̾��>��>��M��%��g4�Yܱ��¾���>�Z��ߎ=3C�>��c�熭�e�}��ø>�b���vĽ� #�=l�>�\ǽ��<���>�.�>&p.�k3��$#Y>�ǽ?oK���9�f*�3�����y⎾ �h>3�	<5�R>򀘼DE\>�־iYe?�W'?�탾򦜾����U�=����y�=�����?^}6?��+��MC�؏#<2�����>В�>�`�>�nO��H?(/A���
�'U�=�|�ˬB��?��>~SD���"��-��v��)��1�5>���1~?�}-��0?7V?j�6>���vW>?� z?�'��Z���M\=Ѱ�=sn>C.n�D��8�>p�0#�>��>�H����;���a���/?m�B8N1�=�"�/Lq�R�=�� >��.�k\��Z?�<�$��)����>�0��l��	����Ľ�T>Ț��KoG>�Y�>anx�������ˉ
?b�D;�W�=m���Ɵ�����=����3��i[J� ҇>�\z=M�6?`�4?��t?�y�>��潦?�N��3���->����'�>���>_q,<�#�>��v���ڽz�>�sl���e=K��>l���JX�������Λ>�e��
ե=o���>�d>9Ӥ�}_������]R�V� �aǚ����zK>;�v�7%�=p�9?S�=����@�>��"?ș�>-��8郾G!�ۺH?��$=��>�)@>{�־*�i>}7?��/?P��X��>�`�>���>�#?L<̽�k����p�I)*>ͧ��]�Enc>��?�ؾ���>���?oM<>\ɵ��-?�>�0̾ ��;	�*�d�>ǘ�>���� 9?���>��A�
o���=@�)�O�L��fj=��E>��>۹`�������:>�{>����sU�=a�=����}��MB?_ɖ��X;�46��:�5>��_��8'�K��>Uf >ȃ>/W;��9��/���嬾;�>��T��;m����� ?�?��6��J�>W鯽��پ��n=�%">�-�{�����m�?V|�>�M��*Gt>�f>������:�}�>����j����Z��HU>��>��?OY�=�3~���?��0>�<?>�𕾼<>��V?�?De��'?r[?�g>󇛾����uɕ�L�Q�sֶ>�߿�>|A�C[��(��>�Ƭ�냉�
+;�䬼>O6�	8�}3�>�n�=��=��J�;���؝=�>�ͣ�"���i?�!���^��ގ���>��u�P&��T�> �>Ŀ\>Żv�'�&�5!k�
����|��:?cx/�G==�hF���>�p<?���U�Ѽoc<&������]8�<�D?�S>.;U������%=�b�>m
ﾽD���z=B�=}�@�e]��8������=�w>�=��=,�{?&�E?���>Ԕ-?n`=�g�=c�F�������G>[.�����IE?�+���*=�>�ư�O��?N�r>�hq�9&�`�>Hh�u���Y�����>���Y�Ծ�p+>�����pya��)�� �5���?
�2��,�>�����2�����-)?:x����j��Y>?>���k�߾���d�̾#4��ݣ>�oC�$X�=�.�=����m�?Q��>�h�>�&��K��6�u=���=#��u?{�>�4?��>��I��w�>`!�˨I>g����?ҿǽE��>���>���==�P��5����>�9A�)a�=��V?-�;m��>}>������ؼ����>UK���*�%6������)�o�E���q׿��==)pk<t'����^?��&�$\ =ֽ�B�>�"�>!��>�z>K`%?��7?M��>ـ�>�l�Y��=�H�<x)O?%ޚ�i5?�'�>� �>���7<�>9n�>oJ�>΃<= _H�w���V;����)	>���>���a��?�����&M:��KC>t/�>�`a���征����<4h)�pT�<����/޾�Z�>.��>��?4M����9���1?ޑ?��^���F>�=�ċ= kS��(��7�k����>
��=��?CO̽��?�Y꾣�$��rｻW}?,��>�6k�Z˥=�>�=�\6���/�b��PҼ��n�S�ˬC?���j�>�T�>���>� r�5#�>�?��)?��μ�7��8�D�Z�����h��>3f=%���_̜>'{~>t���X����=�>�Ѫ�W�<������#?��Z>/w>X��^��>��>���
wϾp�@?=��> �i��Ռ>U��>�_��s�V�A鑿Z� ?ҧ�����>t���	Ŀ>����峒>�<�op$>o7W=o���g9��gz���/>H�??���ھROJ��R4�Yc��8�P1J�#b�eˋ>����G���l��_���M>b04����s�����>�	����`�mm6�@Z=p\���>��>��T�u�нu/�>F��>��M��V>1�f<�p�>��X�eg�5%Ӿ҂Ծ��3�0�?A����?;r�<�wj��)��5�=g3=�z��@_� b_���>�)���V�=��\>���>�=?�ơ>�:�?JJV?\C���*=.��">�h�۷��۾]>������P���[��p`����>����#?�Q=I�6�'���|P?�����[�������ܾ�>���>s�/?��?>�q��Zg>�}���9�>A޾��?t��>	>׾!*{?�1�>l�������x�WY}>_�.>�g'�Y���|1��-?�sӾ���n��>�V�>NO�>
�3�b,�>�T}?g1�?֨����>�V�u>��>�A>	 ���wt��������E>��B>(��>m�|���c�}�>jI=l����Cf>��V�A?d�N�b�6?׳��O E?�Z�=��>ٮʿ3�>O\w��'�>�F<>�wF>m��=�{=�L ���E��o�>G��=sV�>�${<�+���=����J?��d���(F�� >lݷ�4
]>�J^=�>�D
�K'�� ���� ���"�=�;U���`?�[���_?>�:��?��>�Ɣ>T�����!�8a�����>۴��F�>O U���/=<�'�P�����%��*�����<?��>ec�>8���;e�k{�@��fW��5��<D���a�>J�羶ݾ�����?�������-;+�qߥ�@
?��>:gh?7�7?�|�{D��l������R�	���>�[���E?����>`t��l��>�Т>�%�>�� >�+�=l�>~�>x�?����3���->m{>	�w>H�.��>j��>'�>�y��b?��=�6�>��.�Xj便vȼ���H��`��=5A�=�ү=h'7�n�?�'0>b_z?���>ઉ>��!=F���_%�?���/��?@�q>�����H5?~E-�B�U?pU�>�>}UQ�,D^�>�&�|�b{�S#>+@=��NbZ?X鳾�3T��+M�G6.?R)�n��A)?�%2? ,�=8�Q���>�T
�?��vm�=\t�>]��0a�>Ol=��="eV��c�>,�>ᨡ����w/Ծ �#?�o�;��=�y>m "?F�8�q'C?G�ž�~�>>�>���=�S
��� ?�$?m�(?�K��<�=@�$>10��j�S�H���
`3�)�=�n�����>ƽ����=e���g\��?a.���%>�ִ>�?X��;��ýf�����H>}�uq?���~h��ѥ�P����	L��v3���e��,�>H���^Ǿ�/=?J�<Ñ�b�Ѿ�Gx�	!� )?���$�>z���ݩ����>�˾��ԾJ<q>4�o>��>�A������"�E�i>V���5�)?&�>X���A�ӠѾD�>N~/>"c��x>�>CJɽ\�=�0�)�M=�j>K��I�?e]z��J%��?��?4�aj�>n̓�N�ɾh�=>��`>#��>Zz�>��?��>�p�
>Z5�?=a���e�\����?ş�>�O;�?����?�<�=\�&�)꾰�3��j�>a.�=�q��C��F�?���>��?��y>�᯽wP�=���]�H���������=��h�>O%O�� �� �t?��þ�h�=�5C���?_顾if��ѭ��}?�ܻ>��̾�?6�?���<nE-?�������?T餾�=��4=������>(̍�Y6j������'c>�����=�g!��h>/����=>1~?t����_>�<?薦�/�Ǿ��E=��l>��?��FC�_[r��K�{p�>k��=�=?��k���>Fݗ>�޽\�=\;L?��m?L�>����r��"��h;�v���#`��D�=�L�?��`;��T>*.�?ɒ7>�vN���>�]�>�+?Lk����>��>ڮ�>�$�<rݼ���>j�#���u�R��>ʂ=���="+�>b�~>��G>���L3V�ER�h��=<�=��d��>�{x�NȘ?�	�B�<�*��&@�>���J�U�>
���R>��?���h?"{�>#U�=w$�=����Bp?��:>��?����y�;>���=����⵾����{!?��!?9�	?��>��=A�:�\[?�����?��?\�K>X�.?z8r>��Ⱦ+��Ҙ��ӿ%?C�X�T�"?c�5?�}�6L?6=��?��v>���\-ս��$=�`e?2�J>�^s�	�Ͼ��f�����ݾ��%?��H?�;>I��^(s��28?�)#?��!�q��=�Ӏ>b�>"�V�~m�#K��]�?�(M>�(>�嘽{"?��[>�[=D��?��h��\?q��?�Y>�>��5�B������fG⽽���h-����?�,�����幣���;?[�v�Kx���! ?׍%?_j�>�*�`��>~$>P)���,��A�re�=ho#�u�~��۠>�X�?�Ǥ��S�=r�	>���>;K&>����J�=�^x��DھV��4]u>u�A���?��=7N<o�'�c>t������{J�Ѱ��-
?oj�� ־$w�=-��<�f<����;��B��q&�>�>�a޾�P����>01>���>����>�LԼ��߼6��
��P�<����x�>W�5�a�A?ohG���>OI>�%�6@=V������>�[�ÛϾ�����=<�H?Vӽ�V�O�����?󙾂���h��>�j�?�s�?���Ƹ�>��w�>>l�={��=��0���>`���ʣZ=��1�O*H>_Q�>��4��[:�;o,�1.�?^�����=;s�=�$�A�i>."s�]]�>���3=��h��>�B�����*���ľ|�߽i8�>�P3���b����=h*��Q�>�,G���R?)W�����u�?�p?2h5�bؾ���;>�+����f�p�?G��>\��>����ym�k�>�y�>(����ؿ9hs?BN>`�L�"��~�E���?W�=m�ܾ#\�>���?T�*>���>�hM?�#�?��=TvB�H��H?ɚ:> w�>�I����>���R(p�9V�
�?���?��>F���Z?�W����<�כ�*��?�f��T��Щ�W��?����98�����o�K>���=p����q�>��n>��ؾ�+��i"ž5�w>e���nW�Os>_�?N���
}˾Q��Y�9�������6�=Jls>^��V@ۼ�����_>5��Lg�����>���<8 ?���=Y�d��H�?�o+>}��>��
�.����>��G>1U:�� I�+墳{�>/!
��81�kা.
���>	u??�m��*?i�>�ޢ87�Žs����.�ȍ�����#�L�n; ����f�*��k=`�>A�>�������I�;'��>��5?K6'?�G?�P�>L)>��?`-�>ѡ.��e?��?��>'��>V��<i?Aَ?\x?+FI?.�G?�Ţ=a6���������
��������&������>��?Q���	U>!=<?��:���a�m����8#><��=`���o��n>F籽�Ƭ��?k�*��Y���o���W?�dq>����,*��lx?�J�q����n��>���"�<��k>�l�<X=>�W+?w�(?;�>���>2�>�oa�Q�u>��b>���<Ԭ�=��?�s>�u��r���8?��>����f�	?�C��U-?���?V�?qo>���S>	�>\��.刾_8�����fm��d;��[쾇���n�����>��Ǿi�k�r����s.?�a?���<�b����=O��?�gW=߅�>b�)?�LD>�ZP?t�d=��>�<�];�'V����>5#���<����-�D>���>�!1�o����'>!g���@b��8�xkþ�H"�-5��:�T$���ނ��h9��,� Tt�3�>2>�݆��y����=	���P�,BὯi������d�Q ��]\нj\=>ȃ��*���T>EWA�v��>�~h>�E ���"�_@�=O��ϕ?��?���>?8T�#�B�J�>-�f�	�u��������q�`���g��Pe>K��vpS���>*8>4,�������?�0��B�΄漒�?��f>��?��\?�ŀ>��-?�V�>>�>[�e?�~=>��t�[X�;m�Ľ��>��¾�!�����D��ɩ��΢��^���!����[��>J�L��g�EҦ�b�潂"?�;j�:����е?Z�<?v܊?-O��rP�>����A�S�X�>�A�>Dh>T�����>Ƹ?���7�?Ҷ?�u��܊>8.q��4ÿ ھa�!�V����]2�0�g>k����H>��?5�?W�r��>�=ԇ������-i�����>�ݍ�I�Z�_������>HᾂP������!��_�`4`�ݞ��Κ�����>�n>k'?��,?�����>�k}?��O?�p�:���?g�E?i��E&L>�;9>2�?0��]\�����P^?�b�����	������T.!?�����Q���fH?�P��n�>������>��i�x�?>i���h=��㽡�>V��>�q���>��
?/G�?�ȼ�L���
?G�=HB���[��?�Y��>�3��Y½��f�)==^��=���=��>���=ay�rS���۽�
�>-hp�	�Z��ǟ��T?�0���&����B��̾��>�!�5�g�躊�߿r��&�>�:1>����1xe?��~?��;?�|�=/v�>-T����ھ��u�t}H�3��X��>�2>��=��b>,%��+)Z?S8p>VD?�?Dˇ?�@?��=U ��0�>wD%?����\�>G`�=36W>ז��>'�$>��->~V�>����$C�>��
b��@CB�����y+*�����R3?Xy�>{�?��$>�l?\������>������Y?��?�O�?�M�?�/z��w?�L�>������?��Q�Շ�?�7�>�Vz�h�>ꪚ>{u ��b��?c��(�w�>�ʰ�aRe?{b�>p{�>HM(?����S1����;����>ǹ%?��<?���DY�>t��>.H���>�
?�u��|�h�̾�)þ�����c����=r��žl"��5�?�v�)��Q?��J>'#ս��>>���aK>?0?}��?�]�����K߾?�����
�=�̾hB>�����Kξx���������l��-̒�X��>������\#>�?z;	�<-+>��>�i�?�V����?�c�>�Q���&?�p����S��h����$>2�ۼ�P�Uӭ��ݦ?�����=��=����?�v<��!�������w�;�>K�">6]�> ��ZA����>_*�>Bp��{?߻2?��
?t�W�Hp���A����f��_۾���t>����+���p=X����F׾��ʽ���>˔�?b��B�ݾL�s?h�?��>���>`t=N��>�U6�z�(�mǴ�~!=�yd��V�;i!׾�V�+��>��l?��f?��	�=Z�?�>��=�M#��z"?�[y�
�c�AG���6/?+^5�ý̾"��=��O��mi�&�>����E�j}�>p�>k����ϥ�7��eK�?�*��F�S>$��A ��Rɾf/?���>��½�0�>�+��F ���Y���9>��>L����*����t?8-��] ?B���>�9=��>�(c�٩�=�_> џ�פ���־C?�G>��־|�s���> �\���(��G?��C>Ux>u��=�2?hb1��Q���>?�?W�+?�`J�p钾���>,v9��~���������n?�<GT%>�X����>.hu?�?�;>��0�b���S\�>c��@�=Q�ҿSwľ�>�O��n��fI?
,�?��ڽ�=D>f4Q=R[?����4�>���>�<r>�W���)?O$�>�㐽Z4��Ⱥ��1�<O�&?��>ԆɻY����?5 ����>lt�>&(	?�W=;����i�a�i<��=r[ʾ�B��d�>�+`�<ޠ�8騿�{@>��>�[���~���"?���>��4?�NV��&_����� d4�e�R�C�2�� F���Y�u30�O ��Cƞ=a�g�O�,?�<a?j*�>���<��2>4Q?M$?�G�>��?>��>?^?������3>�����M�=8{�������E�c?�
�>Ub?P�D�bB�=׹���#?�z?�X�>
�$��a,������?[[I��$ԾE���vH��Cp�^e��?(�q�׽��{?H��>{�E��<�"m?N{O�tN>o�����>6�8�۽)�0��>$�O�T՝���M>м?>�ޫ>e��?�i�?%��?A4�>�������>F����|<�^�3>�ڈ��z���8����0���?�?�(�=�q*?d!۾"�,��$���>RV?X�2?��P8�>2��>��<����=a?�>_�*?��c�F�쾼oL�m��?*�7=M�����?\��>щ��u.���C��G?3�d�&|7�c�?��E�H��<��^��_��IT>��?~�U?��C���#�ɨH��V�>�>þ>ψ��2>���L����������n�ܲ5��Ȋ��CügLս�
�����=s��;4��ۮ�>�6�?*�ҽQRR�s޶>��>��ܾ)޾z.(>͞:?�
�X�#>��?�/�?�A����j�b����_>�Fa�W�O�4�˾+v�QO?O�%?���>���>�z?���"�?����<��IN�yۊ�Dp$?Ʉb?a=E+�>��^��*羏)>y�=���>�}�=�~�>@���î4���D���̽@]��Ҿ�D�?>�W�=���>�y�z�=hV�>j��7f>���>�A?9�U��?��rp��>�����*�P]�=~V��&.F>��)�C�Q?�2���<��β��z?�m侩C�>��;�:�>ُξVfE��0�=k0>��?
�>�
����
�ixn�����D���W���? ���j��Rۺ>5��>J��=��.��8M?� )?p�L?R4>�[�>p}v?(L�>��=��@'?�P'>��5=���w�Q=�J�@������?�u/?��f� ���?ׇ#?��Z?�0?�6?<4���L!X�����]?�q�Q,>�΂>yv�0�=x�c���m�e>���3��{�� ��������jR��y�b>
�>����DG��䖾Nd2���@�[.��֩��:m�>	JQ��Ď�T�=h~b?��&�����=��S?��?�m�>��ѾE�B�8�[>���>vJ�>�k���>Rͤ>�9��M�Цl�4��䧊�8�CƼ�>�#??�N�����=�<����G?dM��Vξ.}�>;of>ӵҾ��*������}6<�>ș!�Rp=���>�d�=!7j�u�b�[�>��?~@d?�c�>�*??SH�����ϵ�>%#?M0&?	c��ʜ�?;=��:>@�]>ۏ��z�J=T�t?�/�>��3�޾�*ѽ��f>Y��>ʨI��bh�)9�<+ս��*1?_���X�>(�>.�5?
&�����( Q>H����t�� ���4��V�_�N!>B%y�둄>d����:k>�f`>#�e�#A����>���@��tʾo�4����>Jt��v(Y�pf�f^5=�?�P�>
�?w��>br>K�5��M�=��>�s��Վ=�c�?����ݾp<U$���.?�=H�]��>�O����,�=Nwg?�@�>�R%��v��	�7�D>�z��$�=��?���)���}��M���cս���<<��>j����K��K=���>�
�· �����8�>��/?�]�-�>��=�+���t>�aq�"�Y>܀����%����?!S˽�S��{��\�>P�;��G����^�̾(��(�/�b\<������0�?b��'�[l�1?>W����>�����~�y^?k���JY=2Ӿ����6⼟ ?:��׊�M�Q>�q?����c����˾,�>p��>�y��oz�>���=��>>'U��q� �;?���>��!?~F������=������3?�P�=�����X=�ތ�(�>Ǻ3���>�+�>�� ?a��2_���3P>� �0x�����l!2��B�=?�>L��_��>��>�'?|s
?�`�>��6� 	�5%�u�">�:\��;ܾ�<c�|�>}���"$�yy�Y>2>}[�=���i2u>+��>�>����⾂��bO}=@WA��b�<�$b�m���p�>��>L)a����>�<ѾA�O>I�E���ľ��[=�y>�n��6{>du�=�N�'�A>ZǼ�w9">b�þ���=�$j�)оf��>Y����Ԓ>xL�ʾ�>�?�d�<D�ھPY|��X>��j>
N�P?B�y�/>kV��h�m�]���I����������=k�>E����������%ߟ�Dܲ>��>�����<�QC���>($�>�z�#6�k ��e>�(�=틻�B�>/=L]����k=���>Lf�a�-?�.����վ+��J��>���>����jxU���=/��=dɜ��g/���=y�޾/�0��A>Kx�� ?�j�u#!�G��aʾ"UA>�>��ѽ��i��� >�a�>"�#>����V�sO���>:��{܏=�v�>8�־B1A�ߞ6>���>XQ>e��r�>�_�>͖>��?!�T���>=۲N>���*]<0���rN(>���>љ>�7��Ա�n��<�ha��#>QFt�/�>��u>*��>K�=?�>���9�f�վ��=��M?>`/���0>����M	?�y%>���=�žh?��L?���>�q�<"��^�>��q>�b>���J��>��K?��J��P���}>��>S�>�U��&�����8��M��ň�P�����Ѿ�0�����>���>Ÿ��"?͖���s��pi�>V�6?���>��>cU'�lʘ��s?�>ͱ��T�罞{��r��>Øz=�Z�?���Ӏ�k�>P�>@k����y������d�>]��=ɴ���ݾ�cv�>�bO>,!(�Tψ�'N?u�L?Ƚ>$�{��ח�~!�>d�P��*�>^ھ#[�=�c>.5�>#,9�'�O��E>qP4>���� �ey���(�>�i�>
|��QT>�(B���8�[�;���%���>?��>�=����-D>�<����>���=R��=߇���痼�����2��DX��W�(�%��~ľ��=
?�;�MH��;?>	�=ZR�>c	���a>��S>P�?I���� �>��%>${�>b�>�<'�A��o���6P>��h=�׵=}厾K�M�۪��K��>��>�?0�	����}X�� �ܾt��!�:=Ƣ�=ȸ���>��3=Y<ɼNԴ��8? -�=��I= �K�OB<�d.S�b �R2��ZX�{��>�݆�啾,S�<j�<���>	�E>Z�>��L�1U�?r����>�j�>��>)�;?��޾Q=�L���X���Ž����`]?��ֽ�_��:���V���(I>�>	$ܽ�4�=�Fe?��Mw�,A����?��~>+9�=���:犾�A�>����F�>M0��楼~:M��OϾ�($<į輺ʸ��SC>;#���S�\>#�Ⱦ���>5�侇�6�v*����>�J0<���>���>�H�=�����r>�>;����&�˿����??�Sv<0�=s���܏>D�=?=r�8qE�>��^>WK3?�U:�����D=>��=��u�� ���9ꬽјg>BU�rW>'Z��ո=�h�>���ǿ)��> �>utн%:���w�oxO>�u>ĲY�G���H���2�7X�>w�e;�ež�WA!?`Y7�N���y�>J>��p���=��ƽ�D��q;���Eh��(������I�>%�Y>Aֺ>.M]��u�>i�?^iüSr`���>�K?9f�>6���S����>�I*=ޢ˾�*=G�X���Q��&>�=I{e�h�<ij�/P��H�>W�-�_�b=mʾ���@�+�@�>/rP=(��>��?2��>㬴��rp�Y��>uXx�YyJ=��;Z�>Y1;>��)=�E����>���=Y����j7=�s?�Y�<
桾��9���	���o�q\u=��b=@��<9B�=]�/>�	��� ?i�g?*��>ws�>���>���H�>=������>a��>������b��H�>����
>��nZ?����齟�Ҿ����;>��>b�o�ȝh�/%�vm�������@�=-���$�#�J�a�Oc�K�R=*&.�Y�l>��L>�k�����<�~?�D�=Tg���xE���>�>�b���C�=��k���¼���@#�<�)~��=/�
��ѳ3?�w>0ﳾ���Y�k�J�>�٘=g?����u��Iaɽޗ���>��=��������3�>٫�=��^��t�!�?�.?��>�����|�?��>*�н�D����?�r:M��In���~=��>FP1�����y�>�C����
�k=S��8���?�4���ѵ>�����V =�Q4=��>�L��J{�)s�=9a>�A�V�Ϣ��l��=���=w=ؾm|h=��S�֪.��~̾^	������>�>t�پﱼ���_">K��>^0>2h1�\A?3�T� �)���r>�����P�� [���>�N���v��9�>ơ�>n��=����Q�u��R�>n7;K��=�+�>�WѾ(ȼ�6���c�>�Ƃ?ґ�> ��j�r����>���>�9����>e�>�v�>c��>n��1P�T(�=�/�>t���m`��=;͖>u��7�:�Ӿ�S>fMX>*ލ�U�9>@z�>ۺ>���H=E����aA?.+9��y(��4>:�:>��޾���(ؾ���=\>�Z+��ʵ=�b@�����h�>�v�{���l���1>�`v=�u���¾��νdP]�?� ����=Ql��G2?�qK>4`ؾ��X���H>���>��8���*���s<�{�>�8��"�h�a��Q�>��>cU �ř=?t>=O�>�4�=���=R�>�2���q>�F�>B���<ʱJ>Q�R�XF���žR4�>n�?OU��ۺپ�(K��3?�[�=`\���@�v�3?��m��Y���i��z�>c�������	�kA�U���AD� ���0�>�2=7�a���z>ضT>���پ{���.��>��a���ߟ�}�d���m����=�>��=[̹�ϭ���R�>`�f=�U�ݭ$����?� ?�L�>��=��}�>�A>]��=1�?��>�d�={V��kZ�;�׾$�ؽ>
.����V�-���!q�>��>L?�=�[{��7�>�y�>�iƾG��A���=�C>�FǾ+��	/�>,��/P<������=��>
�e���v?��4>�@+?�|�>P��<ן�>hS��v:@?`�\>�O=*�>��>}zZ�0஽�m0>�o'>��>s�U���>轥>ʈ2���@>���>���>��>nEǾ�����W���0B>r��=��S��Sm>m��>�**���
>�?¾��4>ˣ>W�WVk���??����۾/fؽ=����m�=�-?\�>Ru_>-A�<n�A�XwR=��x����=LS�>�$?x�ȾG��� �ھ\?���=:?��V;�"?��>��W��>�o��y�������L>�Ȭ=X%>'f��0q>t�Y>�����ӼWդ>�cX=��>�!�>�-�=*B%��TI>9�?j��>�ߛ=k�Ҿ�b����K�!�
� ���ꉾJ��+�>^���������dh��<��۾Vl�6|6?��]>1���"�9�iʢ>���E���ÿ  �>puپ�>��b�����>ђ>���<# ���?�
?����H3�Y�=��q��#c?�,޽x1g�Ik�>���=��/�U�^=����_��̓�=1R�Fs>׊��?T��|�H�e��[�=s�����0���>�I���^@�O2e<b�i���]?�J�=�{����ľ{������?�2?r� ��]�>X�=�t�ʸ(>�K<���>�D�>DdN�t쑾��%�T�N�Ag>�X>�FV>�cP>���>GN9��	>������=bڐ=��*�znx=��?��7�iP�=�AD>��&>(�5>�r���?E�=�ּ��?YO=���<?�;�۾�����l=�؝�y��l�?��T>Q���S�׼�2�>Ԏ��"��n+??�E��8��q�)���+�>�%7>�Q?H�I?�I����?�K���y�����05���B���˾z����8>C%�>�0�q�>�����b�0�����Ӿ)�>Z��=!g?���\,1? �C<RѲ>u�6��
���&�?׎�>?EM��?�9X�(=��n=���<}��
��>�X�L)�|�>�7*�F���?8>�k���>��5?2㩾�X=վ�Z�C=��>4��~�>=l����ڽ<lY?w�m��rоb�?_n�<�u�e�ʽ�b�+	h>cJ�<�.��)Ͼ�K;�Н�.�(��/ɾ���S�j>0R?��N&���->�uսxO�>Iؾ���>�6���y�1��Ga��W���3�>1�?Q;��%��� ?�J���믾�b ���G�r9�=6�9�ʽ� ><�8?���>�N��?�[��-�=�&�<��#�d��>�	>M#�ظb��.��Y�>���>s#P�Ġ���$�d��=#�������S1?���72��A7����
>��>���>Z?�xa?xؾ�����פ��'�uo��'=�Ac�wj�>/3�������=?��ɽ����C?7�>d�������%m>��>���ל�����>��"�:�>�W�'U!���>8�>�f���<�)�>�˗>�x�<�V�`b>3߮�C�U�SG�?�귾���>�?.x��s�>��?c�>� �>��>�����=YΥ��?nyB<u%��e?�H�����A��>� V�G]?\˼>;����D��)�t�پ�E���9&>��>�7h!�*}!>b���Q?'&
�������>���<�^���+>ofE>�]=1ih>��/=i��ڒ�>�aĽ�d�W�=k;�x�>���\W����=he ?^1�:�@d=���=��'=�<�>��;>�TH���'?��>�G�h�N��}�>QI	??z���=?˫�E�˽E��<վ�/����f�/�*����3�����>L���+U>������=��¾���-U�����>��>!*Ƚ\�C>�~��1�w>["$>��¾FV=>��>d�P?�@�>�lS��khݾ�	����q�>�>�����)��C���k`�+���52=~����E�a�:�s|�>T�i=)t˼��#?�J�>&h�󖿀z>��׾B
>�6��&����7?�����@>�q=�B�<h'���RS<i	žO9�>�jk��hh=ׄ�=]#?��:�|s�>1b�>�YZ�N�μ���:�a�ӦϽ��{�d�����B�>�1���ɢ>ep�>�t=��E�X�l�u�c>��gӆ=�4���s�='�?5�p��Pپ�"H?3�D>��=�NQ��y��F>��*>k�$�����.c���2Ǿ�p��Z���D>���>�?B�`9��}���$-��?j\>�?��?A,��ۓ=��T=yP?뇒>G����e>��C��Ž����<8��=�E?*�>A5=dż[e�>�"�>xUԾ&8,=�W����>��+>�+ƾ���c?\�����Q���f�ھ���>�1?�i>	\��ɤ>���>��پ� ����>�R�� �������g��u׾���>o�>��<��4�?�#�>J�־MѢ�?yG?Z4%��@������}������t��E��W�����>o��>H�0>����_>�Y	��,?������t�:?��
?�X���=tV?p��>))ǾH>���>dv��}u��-�7������þ�9 ��m�=+!�>���N�O�9N����9����U=��=���>hs�>��f=gžǤ����?�A7��-�c�o>@rL��u>��*�a�>jn�>�^I�z� �vPx<dMe��0�=t�:�����>�>3�Ι>N쬾��b��D?_~�>L�>�A?<q�>�@?���=.cH?�� >.����?��7?$P�<e1;�񍢽����ɱ���x�>~�+�x̊?��==/>S�?��ؾ �?�,<g맾Ѯn�h�M>��Q>���tu���r�Fߙ�>K-��-9����R'�>7]�>�B?^s9>������a�>�չ��<�=6Q?Ӽ�>dS�������׾X1?�T��b�?�r�=EuO>��?<s�=��>���Hd� j"?>!���
\>���=�S���;f
�)������=u
;>S����|f�<��u��:M?�?��H���>��=ۋ���e>t�->��=�qν��ƾ�������z�(��w�?#�=�'���=A
W>����=��������[�`������q>$��X��2�>,�<$���	��=s�B�t�.?�B<>�O׾��K^?A9r�3���!/�#�K;Z?�PYe>\,�bL���s?Љ�I�K�i>�!�=���K==��G��J>�I½��a��I�����L
���>��ژ��2?����L�y�O�D>��>�qþ��1�Ǽ�G>�+���E̾��־��=�6<>��~?�������=E�?��>�i��#�>�,>�w?~�
�پ�4�>���=Q[�>�Cd�h���/w�>=_7�T��A��=p�l���?()�=0ƾ�6����>�ic�[$1�'j��1�|>�%n�2�4���>npF>8�f���c=�eF�Pֵ>闂>Gg�t�P�u�&??���X���Z]�o>����?>W!�	�F>~Y��־�Ӌ���*?��ɾ�T'�l��>4p�=h��>M�0����>!�?i �H��8�I�2>��h������ľ��"?�ܾP^t�AU۾��>�>P&��hr>̝�>[�o?�T7>�HP?�-?E�r=j,?A9�>��?F�>�V|�W_��a�!>����� ��E�>� ?�H콵�� o�=�m%?���Q��>?RF�#��>�<�>*)/����2�=?@�}����f�!����>kLS��޽��Q���^>/J����=��j��kѽi��>�|+����K�?m�����r����<�+7��4���Rw������?�}Ⱦ@H1>~��=s�<=o�=�>�&�>��	?i=���1�轗'O?F�5���H?�$0>Q ��.1>��?�Tv�O�W��5���fD�$Uu��S�V?>��>H��=�t?C����y>���=C�4��֑����Q�DҾ���.�#���=O3������)C��'�>�N>$�x>52>ɓ��0?�}Z>xB�>� ?���>�U�>>k��>�X�����?�. �2�?%��>���<Ź��2ܳ>���>��l?�QU>\��>�>�׆����?����Ѿ�F���虭=�r�?��=J�A?A{h>Ug���޺��������H>�=�Y����>�rU��䑺Lk�D���U�>�!K>�p�=�O$��;ս��>a��>�ld�Uq3�~ٶ��>�P�Ο��e��9p�(��=�!�?Nd >��V?�s> ��;���>��+�Da�יǾ���>`A˾JSt>�V��7nz=_~��]1�>,x=[�>�+�9l�=`�!?ɿ?Ղ�>��W=��>��?�Y�N�a&�)�Ⱦo潲�"�ʕ�f��I#= �M>7�Z��㓾�,�<��>�r�-*���*M��n?|�?n>(���cR>H�ƾ�Ǭ�"�=��>�a��U�Ҿ����Bڳ>M��M+� �����>5W�>L������P��=oX��Z'=����� �{<���G��>��ϼ�X�G��;��<�te���>��N|���t��D�NL����;h:�Rl���#�R�v�2�p�g����Ծ	�7���
?�'F>�u�>̉,�Q�(�sW��K�>Pv��،��`?�I>w��>������=�ބ�Ҹ�����\��=�SW��� �fҲ��/?^if�+��>xMK>�Ч��3�܅��v	>��� �=��r�O?+�r��# >01^�+l>d�J?]�>�x�>/bz>��P�M�>�¾�z�=:���
������!�(k�h]��^��n׾T9�=R�
�A�Q?' ;������h�5>.
����KB�>��a>ra?L(ҽ/�<>sz>ީ9?t��=�����:?�W���z.��<]>�����C��e�>f-����
�s�>�`'�)���C��=홾���<�H�>�`&<>�#���>7��>���>�j���E=�aM���>|;��d}��bP<���>|a:����>\����e���+�J�g�	U<?D�������~f2��Ì>��.�1)h;9��o&�>�h<?��Z*�>�_����>8��>3����߾eK>r�?q팾��3�ћ���U9?���=0m�������9>���<�{?L�ξ\��Ѫ�>�G�=���=����^> ��>
3>����[^t>�"�=�!�<�����t�1�Ѿ!�>���>!�"?��p�
=?e4�?�c����׽<��N��t0d<Y�I>|#�>�����6>0�(��L<v�?(2
���"�;eit>|w羲�[>�	I�1�D?�N��lŋ�����A�̵���v�>�-Ⱦl4�M�0���U>��<M�徶m�>���>�jg?�̸>/ƿ>��[=�ۀ����K־�b־�a����>>����>n='>�,�>qe>;�$��K?IY5?�Dg?+�V>�ྍR�>�H�>�Mo�=�P����>A�>c�r>������ >I��> �?����\s�Dk���`0?��'>�1"�6z�e7Z�����
>��=�.�>��?M�?�Ì=<!(?�I����>�.?`��>�ah?ǭ�>��z?Ͱo��/��$?�b}>I� ?�b���{������Խ1����o�+�E�Zݾc��<��f�+'u>��#�Gak=��
?q����L�=h	��Ԟ>�r�>ch?�m��jy?W�ɽ:�>тk��o�>�p��>)i&�wP���&4>6�>:.۽�闾�� ���L?��z��Et>�����L>�)������삾_�#=��J?4�=]��7N:=�L?Ԯ�����V�?�x�>�@��������eۓ���վA���P�=WXĽLTH����=�d,���y?�_�97?^}��S�?�� >)�
?@�	�e��>"S?�ʷ=&�/��c��J�����W=���'V>"˹>��i��;J��o�=>?庾�-��&�o٤�>�0|�d>>��s>2�=�)�>�H|���Y=ľ�>�o.?3z����>�㉽[x�:�1G���F�s=����g�=�m�>�a�>�&���>#���M��?��J���_>
�"o>ӷ>r�{��(?��U>P�H=J>W@��(�2�U[������¾�g��+E/���;�s��>�p >-9��0�>�L%?7�%=�D���N��1�??>��z>v�ƾ�A�>.�C�J��=���v>�1=�棬<���d��>+8.��@�>��'�U#I�s���\;�s�ܽ�����0�LdԽ>>�u�>�_>yu�>��t��=�=Sd�!R>�8�<�3���e�>6*�>�/��ph�t�.>�t��@>G�_?�y^�W.�>z�*<�ϫ����i��i*g������=fZD�1�?�T�����=�����<)?���>h�<[Ub�E�<r���׉>��:pJ=�	�ǽ���:/��>9���!5�
�̾6'�=�,W?u�Y>Ğ|=>>uh�1��>+��>%��^��>G�
?#�@�D�1qo�<|��r�1��Ȩ�w-J���>�V?2᯽�Ë���?�k�>���>����E����>��>��ždK�>�o���o>��>ɤ>N�6�w�>F���}=�O>�*>�i�2�g�g짾���A6I�D��C࿾K+|=c�=�ʋ>Z�X��Y^?�a�<6F�����t��`f���0:��c�>k?*��;?��ܾN��=Gx�=�FJ�R%�>"�����>�Y?p˟�o��\q"���2���q� �i>?���D?b�!��y?8��=T�0���=F�?�����$?�W�>�?o��>��=ؾZ.���B>�<0 ?:�>������>�n��>�b�Q@���=�'?�ٹ�z>s���h�=;�u>C2�֒v�X)��B��p켧��'/v>���=�ҽ=N�ʾ�C=�j�>^��>��*������2=[v?0oP�w⺾P|˽U�����=�a=?5G񽡟����	?�N>��7?}��<�H/=&�>�� =��˽{� �(�v=|D羻�����H�.5�K�h>7KL��<���>����`�=��_��>w3�>W^?�X�Y�z?�أ��Ġ>6w�>z����>Z�7�Ǔ��J�>��[>La>��!��>�>�J��>V�/���>��+�v&Ǽ�ߦ=�v>� U��}>�y�;��zS�=�Z󽛛�>GȾ�Ҿ�S��@�>�ڀ����*��'�t�^�TꉾZ���P����p�ힿ�Ū5?�v���>��U���>�L�=��9?�7-��?��>Lƾ�$>)�o�^=ϼ�=�AF>E�6�������e?�9=��>�wc���>����#\3>S>�=��J=�7�<�s��y��B�=nt�>�	>�.*�uŏ?�o��n>��9�HF� ?���>����>�]5��5&>���U�վ��:=k����>U璾���6��)"P=\��<�z=,-��LV�<WZ�>\�i���L>���>^�����?>zv��(7Z>����ձ��b�:���*>l@V�[�=�%�|�B��ۆ>�g��^?��(��n-�ne?�=���.�s����`�wz�>A?��ҾI�J>�G
>�d ���q��/�:1>X��=>���k�G�.\T�-�>(F�+�D�jw��q��>]ؾ�3>T�ؾ<K�>��?k��>O��>*>*���M���Ⱦ��>j�;�,齏ʘ>ؠ�����b``>z���4�>�R�f0;��Q>-�>m�#�)v��G�о�%?�x>\�2>Ҩ���E��aK�c�H�J ׾@#<<�(�Χ2�>�g>�۠>�6c�*Qx���0��'>�O��5>����1?��=�!�A)��4��'w�ƫ)�7@�"�;�˶���b����>.<?��A>��޾%��Ǵ�s��>�>ɋ佢<����?P�A>;9*>��]>9��d��>&rE�?�Y�����O>�	`�aۻ��]s<�ڛ>??�a �>r�/�^�+>��>ل>B�����оϧ>����������z��=��&�M��Dľ�`D>�Ƅ>ii��L_�>:ν>�]Խh�x��>y]k=�����>':�=,�<|Wl;��=�La>�z��ƍ=`4>�| >db���H>��>�.ս�<>���>)6H>�<>:Q��L�}wA�*�ھ��q>s���������>xa�<�蔾�炽�x�Ƴ=J5}�Zk�� 7>c�[��ҥ�v����;7���?�6�ػ۪d=��>B`.�
���!��a�M>]3��en��h>j�>���ra�eL��XQ>�6>*�2����8�>轛���i�:2�>�S�<:�ٽ�����r`>�� �<��y�������ۨ���!�8�=�t�<	k7�.��>��=��H�IYd>.I>�ca>+)h�G�$����%�*�(��&�>����Y	j��s��wZ�>k`���ɽH�g�Ƶ�>�q�=��=��L�=(��>i�>����#��	��>8�Ͼ@�'�U7�<��m>ɻ�;s5��/��R��>ս6�,����:�sӱ>���>�o(>P��K2�=Ɛ�)׼^�^�0��|�>��Y>@��_�=�
��h���iൽ5w>��E�=���K�>+�.�*l�=Yl>�w�>����
Ľ��Ⱦ#�>�ܽ*�K��C�<�k?�?r>9��S���X�*��.�>�:�=R��$I�=�_׼sw�=���<�J���=��>[��;!����þ�ʾ��	�=�鮾����Ȑ>1�=[V��@����[.�r�=�Gн�����>��=���=E��d��P>���!½A�>�[q�����C�=�2J���	��;�����:��4�=u|ἣ.�=��<���>Vib�26�]��=dT <}P���/�r˨=d��<<����ʾ��=;�c>�Κ>%�q>d�>w���*�*T
>� ;owy����=xU�ȟ��ܒ��T<y=6�n=N��<5=m��[�<��ս�6��S���?+�[;�+����A� �󫶽P9�>Ԏ}�5��>��>G�=�c��Ղ������>�;��Ӳ>���=Ҳ4� ����;�8$w��	�=1���qK���>9X>f#��+.��p׽Nލ>"�w�M�I�`>r�1��6
>���>,,�>�1��=�}�=% > �p���;!�S�q�A�x!^�:��=]_�;x��u�=7*��;���@p=���>^�C��������f�>.�*;V� >� e>$>+����#��s=�n.�&'����>;�>ǁ���iX��*>�����b�
󦼸�<��#=]P���;�[��>6�=�#���RԼUa>��I>:n�=S������=r/l>�6m�b�R�L蒾Xw׽8nӽM��>�o"�9�����=XU�<��J��ƽV)�=�*=@-�2����>%Q>X�>[�">�8S>@� ��8U�z�d�v�s�熒>��c>��m<�u^>�H�=R��=���>|>'�ݽ3�<~x����q�˾��*?�؁��.�뾞��)�=�^�=}�?U�p?�;�TI>���b&�Oa)���
>�>�e0���=��н�����?{ߧ�V\�I"�>!�U=}��8�?>�Q(> %>���<^=ù�>������+>�=/��=Y�<����U#����>�����.�= bŽ(���ΐ�O#���2���	�=��e�W/?�A�=܎��ZTQ����=�U|>g�>� X��uC=ݰ
>2ս��>�UU���O=��=��E>��辺���s>kR>p���r�����c�)}4>jo���	���h>o+N>r�B>[�1�k����X=�VK=f�~>�!� ��=�A>"�=���#o>�>���X������<Pj�,�۽�^������|Z>�t�=C����<0��>6B�=N�+� �̽&g�=<�=�V_�E�M<H2X=
��=0=�>^=�kR���ռ�?i���� =LA�>2X��'׾��o��G�=�]��^��.=tD�>���P�=\�>.����)*>P2P>��ؽ�UG���>�2,>�R�=n'�nҙ=�XJ><��t���1���*>�6->,0
�v[!=���>cI�������Й�}�c=��D<QE�&n<�E�=��q=t>�P�~E�����=�?1�þ�,��i>���v�v����=l����k�a�-=�H=�꠻��žî>�F�� �
z+<�T=��=b��=/����>��~�����E�~��qu>lR�>�ռߣ��x���˻D��=\�}�^�:���=��<��Y��D<~>$>{5,�C�,���;��P��ҳ��IG�>�t=�=�1��>�� :�t��*��}�>�v��Ɔ���q���>�|=�o'=ޭ�:`>��%>K���%? �f�>!\���������b�4����=�R)�	���wp>��p=�4�;3^�ͣ��Qc쾵�>'��>�a>a���3>���=�I��#j��������Јo�$i��H��"U�<�0�h�ʽ����,�>-�꽙A$>�>�l��	��%>F��<W�8��\�������C��{�'Ou��դ�Ԏ�>�����^����A�>(�<:�$;���>����Xԕ=.hU>���=���%f2��h|=��m>���
lZ;sY�<���`�d�@��<=���IJ3=�'�=�P!���t=�^��������z��)�=v�~� ��0b>[�=Kݗ������>�*'���ǽ�=�3�=�0r=C#=�눽o6>C�>�"��ս�b��\3�<�̢���!�X�|�r�����_�¿N��A�/X>�9>���=�ԇ>��>�{��V�?S�>�̅<�Z@=B}>"����9�bF'=�)�=w��=��0>��5<��N=�龧/���IQ=���>0*0>7�@�S>�y >� ��g�>��>�贾�潐xc������E�ێ��Xq$�@>�v.<�$�>�uJ��#��������>�\X��:ѽ��=�\>[{�i�s��T�=m�>_�)�C�>Wz�=Ш�=���#j>=I�>�T��G�>�D�>���<KJ=���؝������]G��$� �:�?>�$<�v��W���P>�I�>Ef�>��G��> ��=y�)�_�'��@-�u��=!�.<��3�l>Nm.>������=r�]>�<o>�ٽ%I��l�=� �>&Y��-���B;��>ý����n�d>6_���=���>ODP>�\��� 5��s��SN6>wܽ'��~t=�;>F+�=�^��뫗��8]���>��<>���:%�=���>[���B�]=��xSN��Ӣ=?&��Tݽrt=Rb�$�>�+ɽ��c>��=L߾B�=�+�>�o:>���m�����=z>����7=��V<���=��r=^��f4�>�ɽ=�x6<sSU�G�<��>)c�>4u����=b8>��|�����cڥ�v<��?=չR>,���?7���>��E>ͽ_2o�`�����k>y���&	�� >�W>0>��Ѽ������}>Z��;��< �>[;M>gV�׮�MsǾ��>@*�d��D�<��>~M����ƽ��Tp��hI>�鋾��g>�_3�m���t�Eh?z�f�̞��>yه>j{5��#��k�t=͘>jar>Z!پ|#�G��=x�d>yi��?@��8�S�t>�۽�#H�#]�=s��>	q�>�Լ�N�;wa/?e{��1kE�i��>n@\�	b��j2�>��g��+�=���=��m�ƊƼ�k>�}Z=�_v>�:����>����D8>���=��=���=8B>�+h�>�9�H@��yư���S>���=����-xɾiO�>�Hݾ̢>[#>��>.��4�0<������>@�������s��� ��>%Z�=�Uý��~��Ց�䂾2��=��k�	�>0-�=�mK��~��>�|_>ߏj>>�*���>���>�����'=�k�>*1P>"�(�a(c>*��&1�M�L<��>�FT�#���g�o<y�w>��:�.��Z(>C�>Jʔ��t��ZC���.���g�P��N���E�>K�ݽԾ���_>�!Ծ;�l�:p�#����>A��>���>���>���>f�/?Tv�>�&�>c%n>!��=
Й=��=f%L=��%?���>���>��>�a�>Í?���>an�=�7�>r�7>�>�.��?d?���<�>�ק<Ҁl>D7�#˾��۾_䰾؀��J�%�j��TO�.��ĐC>i͘�T���Ȅ>�9��.¤�s� >�tž�v�>�P�'߾����|=�0�JY>�>�P?�B��+Um��sF>6]�>�37��f�>�c ��`�>{����?'[0?.��?�y��?_ݾ>��'>Z�#��^�
z"? ��;и���*�>�Û�X}?b�=���>l�=?:���""�o'�=�L�>]٪=Yz�P����>֊t=*)�s�>��%��ƾē�G���V�;L�]�z��=�'����^+=�g�>T��>�r��j� ��zB>��V?6e�4k>�j0��;,}�Wց��޸�HL�V�Gt����V>��?�Γ=��Ǿ����=�6i=��u
�'|��	؎����]�>b����:>��S&ž�%��V	�����Ę��F�D�l��c>���
0'��9¿���w	�9f�R �������<?�u����9��$�J��>8�a�=d>r�m>��5�t>/A>�.��c��x����8?1�	�V4龤4>m�>@H
�F�E�����ھ2)��@I�s�b�t�4�C�o>5#Z��o�"s���Y>QG���0� ���J+�FA@>E��E�8��)?}��G�%?���=�d/?��=�f��E>���?`�ü�b*�]��_�>���>���<��ܾ�<B?B>QHj�c
�,(?�&�=]�r��9&�>��==?������x���H?hG�>.��L[�k�'?��p)?7w�=h>hz��z*��dIr��>��[4=~��	C��u��}2����;�oC�(04���E��>�>ۧ,�{�)��Q
>2[�>�K$�J6q?%��>�#?����uʯ>#���]��u�5Ϳ�ŉ��z���Z��BA��4��vd?�_��l"]>w��=��?�a�>JD>��ʼ�g?1�1?Ժ�?��	?����K�~?j��=�8?Ľ0�f茽qv&>mz?��K�SRl����Ǚ>�۾��^>��t�6?>ai>c��>�ԭ=��L��ɒ>z� ��L�����?��1>S�>���=�������>u ��D����?7F)����>�.B�/��;A%�=0�^>���|l�\L{���9?���\?ީ�?�(2?�����N ?�	>4��>!{\��=��������>�,�΀��f�<X��>��P��=�>a,Ӿ�����1T>�V]�#L�o �=ѠE?�#����Ǿ���(��>�S�>X^,�s�?�?#c�[61?���><} ?�mS?�=?fa�>%q@?��?�xC>���=j�^>H\_=�j�?dX��
��΄��RV1?���?3�����>)�?+8?�����?�g�>5`�>�t<���>�S�>��K��>��21>w@�>�Lb>�o�>5͇?qw�=� ?�~�?{��?���s��>2"%>��>2p��������� �����P�����x��N>!?f�$���>Ly5?Zd�>G ?�9>�ے�Z�~��^�=�>�	6?S�?��߽T��?`8?^!?)oX?�<4>ϭd?N��>s+��������<�Y�>��m���G�(�(�HD�S3ƾ�߾9M�;�H)��]�֛��`C���/��X��I$�[��������l��z�ʾG�����pZ;�f���꾾@2�=�֮>��V>�����>:[�>�f���&��K�w績5!W�ф�=��_>���>WҾ���>ϰJ?}u?� >�ͧ>���=vf?X�c���F����>|��>7��?���N�\�"��i�>_����'�y�3'�?s�I>
������g?@�;C��%�g��b�� ]�>�ʾ�8�@ ���#��Ӌ>"jf>k�.�	y�=$ۏ�(���?�>�k[=�Q�<6�������=�z���G&��5J����X;Uv��	A<��H�3P��O�I���!'���n��)��b��C\�����O���)��a��hȾJ�Ѿ<0��a.(�4dV�l\g>ވ���R?Y�T>�����!��|=�9�0���⌿"G�������ط����>��Y>�����}��{Q��O��\�=7�y8������C��!W�=R���;�=�D�>������U!>��7>�i��P�?�?[?��T?�/`?:�(�:V̽����q&>2��5�Z���`�Cw�ľǎW�tޕ�>�>sB���:(��'x���>�f�퇨�=�����?%�򽲾���QZ��H��طԾ`�D�=f�&��>�C����>5,>3??_��� �=֢=�߅�ְR��4�<��Ľ�m��2>��پ ��-����>�b�Y�}>��>��z�=5��I��7��K�׾�r�����>/#ּ~|
��~9>e`|=��=���Ѽ,��>��O?�k�?%���zC?c�>��?1�.�vgs?�+`?Д�>�r�=�F�>̱^?���<��F���w��� �:�.�Z��ç�����/�c>ݤ;@�����g>�g?K�x=~.�>�y�&�-��s���F���Q�=��w?�uR�!���n���P>g�����81f�F�B?��Z�^�`<�����>>cT�hn�Fh��]4>
�����=� �S�6?�ｾ�==E�������l>�<(��?�|�?3��?�?�E??K�S?�Ma?{�>��s>è����->D�b�3�����a���<��u>9���=�N>C<�>؏¾h��@���9M�>Ȗ��C^��q�S���?"D+>�*��J�5�h�Ӿ��*�">͎�>�l�>��>������>Zmb?n?�(��10���-k>.�j>=�0?��6?� ?��>�ԣ�I��@�=ـz���߾���=E�8?�z;���~�V�=���>&�?�N�T�>���?�&վV�>+?�(A?�#?[>6�?��5?��3?Q�>TX=ॽ>�f�>�:G�4�>�I_>tȈ>gm�>�L�=ȣn=s��d�P���>_��>��f>�t>Nn?|�?<~�f\;>�E=�h�=L�	��*޾Y8���/�9	����	��������f�����6��;Q3���[���䎽n��=ݶ���]�R&'�Ҝ`��C>;}�&>�|����F����>R�����0���?�o��W�=s���q���C>�;�=F�0����> �U�?�[?U?T��>�s�?����|X>S(�>��>�1��i�=!�����>�����=�Xo>ph?r�r>���|H=�f� <U�?�鏾F��>��?
G����>]?̥4>M�p�\.���� �6ݾi^b�*Z����'�>`����ּ�Tξ��־N�=�^=U���+�4��߇�������>�.��Ԃ����0ɽa�� z�T��Um6�f$���>��>��ھ,���Қ�����P�^?�F[�9{!��!>�f��pfD����� ����r�m>y���a=��W1�����g�G�G�>��(��������"?��<�� �]"ƽE�=:/��7<�',6�e?N�?�Na?)?��6?�Vv>�ʀ�����>t�ﾽ:�P��=��>SL8���������k?�Ҁ?z�>[�h>�Ie?ғ�>
������a�K<�@��k�V��*�>*Y�v
�M��=�,����>�o�<��sp���-�f����r�������)=P/���卾#�k�����B�F[+�*U�%+�=�?�5���1�禾���<���>h�<�0���Z�=7�Ǿ�M��sE>.W̾ �.=Pl�=pv�>[;�>�m�>� ���>��мTdb��k�*�V=���=lZ�=��$����=�c?��+��>'�=�nϽY%>l��>/sN���p=��)���o>�^i�+�.�H����� ���'�����'s*��֏>G��>rR>�\�>"N>���>��>���>o�z�݆n>�4�<�S?��>��m�%oݽO�>��A�>��X>O(G��i>�w�>���>�6ؽʼ���詼L>W{l��d��q��{_H�	W��j��>3�=��)>5�>E�p=��#��ʼ=pL���a��a��/��.?�=����@�6=�'�=w��<0��
L>R�>��\>����K�P���u>9��>9����F��;�>q�y>:Y:�T
��X�(��>��> V�>��
?1N�>>oҼ�6�=#>^>Y2>���nI;���ν���>=�6�g�߼D�=�ȃ>��8�p��>�I>󒼾K�A>�P?J+>�������=�\=�d>���eP��]:e�'����a�����>��F�yn���JȾt?��_�bq���#sq?4_=F��n���v�>��I?���="�y;%5?]b��8ﾽ�O��Q�>� �+S�9�Qg�>{�?��!�<�ih�=�>3���̶>��Z=�@�>����%ʾ�f.>$�?)����;�r6���/��>$>��V�F�rS��m������b+?�o��C?�z��� �>�|��P���M�w%?�Ӄ<�4���b��o8v><Ʉ>�,���֮������ ?�Ӧ<W����>P�>Df>u�ѽ�݃�����#�>������흱�`3����I�>R��w�4>�h�>����+�5��J�<=�>{38�q����2>�f�>k(=�Z�>��H>�}>�"V>z�>HF�>m�q��2����=��5=�I�=����J6��ܲ>���<p�S=1����I/>��>�B���<A��>aw�{�
�����a��>���<�
�	�#�̷�>Z>%2p>�B�>��?m��>��>�)����<[�����ʽ:�̽�^��Q@�>��~���ھ-�y>��}�f�w�;��<�5"��[>��>G_�>�Aľ37�>�
?ZO?e��� ���1�>-��=޺��>\gi�z��n<Cŉ>��,�=b"=�&�r��&?3v-���9��n�>6�%>G8�>�F>���<��>1T.���=�\��v����>0��>�S�����.0�=��>�M<:��3u`:�G^=��� ���y�K���׾��!>Fl?-��^8�*��=��>z�$=
�$��3νX��=��=T��>P��>>��>����L5�/m���ܾG��?oJ�;�Qݾ��=e�>��<sZ�<��3���5=���=��&�T/��<��>�;��s���e�>�?���=�,���5��b�>���=�y�wV���ޝ��s�������>h$P����*��>���;`'�^��s�z>6��<��߽��(�ޙ6=�">�G?�R�>��K?�ʏ��>=�����Ο�gi�=�*�>�]��>F�N��>�?�u�>�N�l~��t�>��="�8��$R�9��>�.?Ȫ>X���ھ>�c?��f?�=/�B.h�S�?���>J�r������=9��=W���v�,>M�=2D��7?���=<}=6�?�o>ТG�)��>���	�}>0ċ>t�ĽIb">�>�mM?=�=-uǽ���>�'�=��;�&�>��2���ɸ>Z�$=���>�<>Cl��>�ͩ�j\�>9���������W��>~>�>� >�g���*�>$�?
�>[���y.{�a�I=�==贬>�L���т�t>#$=,�־Qp�����N'>.���c��@����>��>���;�8>��>nL=�|����ȾQD�>9��>&So=MM���Jj�؏>��*>�|�;�w����E��\<�8���;�8�T�v�d��xֿ�;�����>�1��ﳽdvv�����j�=	�v�u��>�^'=Y�{={����<;����>_H�>נ���ǜ=hg��|�>����4+��쥻>7��>���.{^��~�>���=���iD��mB��˝�is���.�=j�پ��:����>� ��.�<8���	?5�Ľ��">�V�����-�w���q�ܾ2��=j},>K'�a'�����+��<�K3>��۽n�=�'=��`��c���<7���8n<pu�>�`��o��Sؓ>r�)�V9߽-��>�����>f�����6$>�J>��>Ֆ��&��W����q>�X��ކ�E^��� ?�V�>���M%>�c=�;����Ĉ0>��<e�h�*�>�8(>�X�&��>��=���#4���{����>n�-�)2��L�=ڋv�v���,C�kÌ>��i>��>�0�>�l�=�ۢ�bn>,��>p���w��\M�=�@�>'�<�QO>�.h��`
?X�>������U>Oq�>NY�=�<b�t�&���<иw>����jؽ��=�m==��R=�)>�&�=%ء�L??�?���>`y¾�q�>��>>>��0��P�b=�>>b�>Dl��6d��eu;����Y^�>w��>n��=��͍�>h>�>
G�/m=A��t�=�/�>���o���0⾽n���B��U�!���8>A�`>)§>G� �.��=_	?R@&?$���󉾮�
?��#>�څ�6�0�#�,>Rn�=� ^=o��>-�=����i�&=jJм�S=Z��!Sݾw >k|׻�l���<�I���9@���5�e�T>O($���0>L��>��ҽƾ6�i�>�d���T�&<D���>f��=�B#=���=�>�œ>�?2��"���>]$	�߸� �U�<�o��>߰�>V��*�e��?�6?���>> �>P%�iG�}w�=�PS?gFʾ钆��RX>�������>��s=�+*�<^6>�!6�'�>�8�'�>�?~/?
P��	�a�>MS>7�>Wq��/ұ����=\'.>_���Vνh�þ��M����<�=�v�>���>0l�>����-�<��>�r�>+y����:��C�>��n>��iY
���T�>���<�5�>s��=��0�iĶ����>~D�>f�:�����+>�+�=��u<�Z�A���&�ès�μ���J>�&<�X�o�v�=N�>��N>�s�=tI��k��>�\�>֕>��5�Z�FE>#r;'+�R��=�=��������?�����U ��8�;)�>�����U����<��!����	΢>��Z��=�>J�%>hp ����0�%[�>ȭ��gk���ڽn�l>��=�8,�6�=����Z5X��=񾢃����=�A�=y����J�#=k~�����>������;R�˽��%�XC�;�������<&(����������Y�>_��{)��N(>#�>����ճ��ʋ>���;\��<�-:�Ů��'�>�(>>n󚻚����>1?�>�Ҿ�;�=��>�=>�ı��2��F�<�C�`\�>=�������$�=�p�=�����<]�~}J�g&y>]S�Ҿ����>w,X>�M�
�,�^n�>�xz=G�>�D6>_�[>Am-�뺼˵�ӯ�>Nq�����-ώ!\>؎=�������5��O���">M ?8ʸ�̾�!�>i��> �8>����b�Z}>a�>L/�ߞ��|V�>8��>?�����9�"'�=��j>�������:Y�jl�>�9��>��p�*��N�>ޤ�>4�6���>��?�]/>�(>w�?��*>�N=�A�>bϼ��7> c�=4fl��ң>b<��2>��M�3>�rG?��>���<K ��5"?��>�򑽲��<>٠�=�'*��*"=wS�k�i�5����!���J?�ؽ� o�,ʾy"?�4<*n��&�y�>#[�<Z��"M�7�>a��Ć��1�1�սt�����F��5�>4q������w���5?�޽��d���ھ��?�v�>�=��3B,���l>XV�gI?���>9��~�=�F?t�1=Eнw�@�<�U>��_U���JM��cp���W�>\��4=��\�Q>��l��������}z>f�!�D	S���ݻ���/�����TM��� �=�B>�>�ӟ>�(>�+�>�KG>�g>�H�?�!?.R?��>�0�>�U>�I>�]?b�Z>�C?�Ƚ���>����u�t��>��>��K?�^?��	?�T>�cڽ[OĽ�6>�v�3>̖��� >�W>��>���(-=4s?7*I���=���������� ���\?�5?�`F��ď=6�>�2�>l�*�_>\
��>�I��u�#����B&"?h�*�~r�{]>Ddk?�R�>�4?��i>�v,?��=���= �U��n�>��>c2'=�=-��?+/	=_Ǿ����b�?^�<?a=q=�|��zi�^��ۿ�=��'>�����S2?���?X��=�>��\�;>����ܪ�t������jL��:�>�>黾F��=���-)����(dW�_�_��?���>�پ!B?�ޙ�_l+���_���j�����>�@_>n>�|�=�#ƾ�
�?x�m�oR>2?��L?3�B�B�@�*��-]���>�W�<L�M�[@����!�Q�~>yP������p[�=1z���\�>�c,�H���Yܾ��-Ū�Y��>�	���Nu���=��;������'�(�^��Y�>�{8���>�F��J���>�����MZ�!�t���=��$�<Y�m�?��;>�9>�~8��i��<xe��.�1>�4>��S�iYU>��^>D�4;�~<�O6?���=�c���k#��Ѽ�Ck8���?~9�=�cJ>(���
>�1�>�(A>�ؤ�>鈽�H�]1��)�<�>�g���>_�׾km�>
-&>���<[��=�v>�_"?�$�>�Q����!�-?I��&k� ̾I�'=�
,>B���(FJ?G~�>L}?�|=>�I<�A�<��N�`�q�=>�>F)־Ԝ>��*���=�>/��b��k���|����\���x?n�>[o�=�{%��3y>�hl=A�s>�F(���?�'?��>��D��> �<����>��}�6���'��V�=�����
�:�¾��=>���$#"�<%�+��u9���]>�F6��a��7��>�H
=�'�-�
�gZ�=
f�=H{]>$�'B�>��Z?��?t�^M�>�?�e���H�i�>O��>^?��$?�~�LZ?pT'=Ix�=���3�$���޽6����o�>�@��5�>5{z?�{о�D>c'�B�A�pD9=Mx�û?��C�<��>���>ي�>%�z��^F>�g%?�I����v]8�"ˋ<���7���6���z�2뾽�'��=�W�>�v�>��#�$O����=_��*�����>��4�=S ?$W�>'�L=��9��N?�ž����A���P�04�>fY>���>�H7?��*��8n���=��4��MX>z�F><�>��>���>�X�=B��=�'1>�tG?3>�`?�@���?�7�>6�d��^��)�>���>z�>�@Ӿ��M�+O�>s�>��=C��?�/�<�?��>H�>��k�V���Ӿ] ��և;��>O�=Eꋾ��J?���i)>��>��X���*?��=2AJ>5,�>a�>¤վX�?��?�ª>*�E?�΁;�t����>-gl�Qk轥#��Е?�i>�G��=Rq?h�>
�yW3?̵\>Hu>oxP�S�=���>PF�>]Ӆ>%M?5�=��>f�3>�#&>n0��r1���T�>��-��-��n>�	g>�1?��"	�_����#o��[��:U�>��?=���=�ݜ�J�ν\�
_�>��=�Tƾ�'����o?�=?��;>�J����<�-g��K���Q	��>�{�=�Fw���+�l��=�y?.�d?^��4�=�j�I�R?nLc��������>�:����Kݾ��Q>++���z��|��$���)>f���4L��n�����=C�4A�=�v"��K>h~���qӾI_�=�뎾!�>|8�����ʈ��k�>犙�R`T>\�%�9m��`��3?9p��T>����(>.H �\�n��*�:�9ƽ����c�6�iE?ie�>}{ �Sć�i>�+����:����ii�=�M7>����ۍ��>=�_u>��G���>�`�>����^��@�")ѾH$�	���b>I�Q���?�*�>a����&�H���Y2?KH<V9�Q'ҽrQ?�@����⾽�h���3��m���"
�;# �r����>&�t�}2�4�2?��Y��i3�OrW�t�Ѿ�[Ǿ�+"����>~u�>�x�>0?�s潊�=���?��I�y*�����$����2���쿾S��>��u?�>�I6��߉���>���>��2��Om��o�>J��<�t�r�]��BӾ� 6�����a-?��>Vy�>xR?�{�=��E>ՆC>\>��S:�V{}>����N�=Ʒ5=�c��o"�df�q=�����>�=Ƭн�{Ǿ��>k�V>����^o?u%�>ҥ�=Ij�#�p�Xlļ��G��=A>.�*�2�?�h?Ⱦ?>d��Y�K?� �>">�,���m�>���>��>
D)>L�?��O��Z�>�67�%��==�徱y����+�_.�=t��>�/�v��>2�����6��>� ����dY�=#�潖ܲ>��>Ŀ��W�*?��J=m��\t��ZM
?ك�;�k#���+�_�t<����}��-(V>�͊=�I�>L�"�cȬ>�Ҕ>��½ō��+� �	��>_����t�����ˎ>չ�>:�>0P��&�?�>S�>@��>x�>:�?u+j��R�>�CȽ�ɾ*�>�g�>��h����?2{��Z���>�r�>W�;���=��h�i�y�E?!> �b㪾t�?��i?�3��Y�^tھ�P�;�����K��7>�?��?d;�>F^E��??�̾^V�>�վ0��=o =�J??��v�u��>Ժ!>e�?@�=a�?A?m�����+�N��2?�A�>��W�r?(?޽J�0?����Ɇ�;��BS>�͇�nnj>�}?v��>���<�c�>��p>N�C>mlj��zF>?�_�>݀�>��T?����p��>��P�6�3��[�>��ݾ46�=��Q?a|>���B:���n�>�Q�=k2�>b��>�v5?(�>;Z�? ���B]��y���'�i�=�ƾ�z����,bE>������O�Q�}��1�j��/Ck<�׾�N��9ؾ�`	�X|���B�
��>����"ϝ=��ؾ��>\�?����l����>���>��T��̋��)�;��=�۾c�u>"�>r��>J�y�$�� =.� ?��;���<ާh?R�J�dXE��=�B�>O�={�Y=��$�B?^�U�{�U>�@��Y_?o|+?p��>��:ɦ�k!����>�CA>Wrz�I��
����<t=���XA�δ�����=\5ս���eJʾ�s��n�@�%��1�Lu�>iL�����~�־H�
�^�ž�莾��g�->�1�<�Ҿ~m�<�	>;��jh"��s��8��i�=$aM?:���iT��~�^�}=�7`>ζ���#��MY >���>-��"�ھ�#�m?=�=(���7���Nl���_�<��(�m����Q���>��Lk��G2ڿx]��͔��n��j��I�?�w�>|�2>�J�>�_?��Vj�>ւ�>��^���?�(�>�����^?}+��nB��R����>�/ռ�B�>F?O�>�6�È��Ȯ�>�w�?��ξ\���{߾�?�i���?�=Ž�Y���]Wn����<�=h����<`���W��ľ5��Uވ�9}.<�$,����>g�F�핾KG�<4�>��=�K=	��>��d��m?�b^i?i�v>�%��"���=������Ö�? l�>9i��?��D�>��/�;��>�n>��I�{���s�羃�[��L'?�MB��?S?��k�?+>k�U>��>I�q�ƈ�=8����j�KU����P>tվ<{�r�>,���qy�Z-�����9$>]c�=DW>:ˍ>��:;(�����>&����=�ڹ>�'?���>ALH>~e,>��z��l>�7+=�>~�>n�y>ks�nk�=�<��_ٽ���>�>gP?�/�=��˾��+� ���<�Y>-^�=?�(�<d5=*����01��u�"�>�X�<S1�;�>_I>52�F�+�(��ES>���;��K>*�>�l�����O^=ž$>�&���>�ȴ>�ŝ>���2��ER���>��=�^0=�'?`�>���=í>P� <�c�&=�k�ɔ�!)�>��o�&����k�w��H�N��	�>�Ψ�S ��'�E.�=��<�_����,�>bBI>P-�>�Q�u����*�(�U��X����<�U���&��t�Ѿ��S=����Ɨ��`��P��=�ȽF��*jO�jFp>G�>�q����Ͼ��m>WS��� ��+��W�=>$S�=��ƽN����论ןk�8~�M[��#�>�w�>v�u>g���T>��<��Ծ��� ���}޼��7�4}]>�@]>SJQ>�����p��3��mi����.qݽ��=����yV=$Y��僧>A$�<�x��`�����T>c���c�� �;�/�>�Z��m�� Ս���8>QJ�<<E�$k��:��=:���н�,TI�Hi�X��>�2?��ؾZP.��	��d��p�����=a�8=�~>x�=r�\>jUսU�|��(�ߦr>�U����4��j�>%�>8w��=�^�=�$�>6�+?֯>]i>�Z�=�I�r�����t�!!��E�����>�)�>T?�=yF �{���=�GԽYc�=�E���u����<Xq�=�z>��=9;�����ɠ>��>��>i��>a��>O����#=��I[l������_=:�=� ��]�>��_>�׽����3@?�>�W��%z��!���ȁ�c`>É�=���>�K	�~%����=�=���o|�>��X?J��=q��Lߦ<ݡ����>�T�>��->Ʉf�͑��m7���Z�(U!==�>�ҥ<a!�=`+�>%���>�WM�P_I�3�4?�Ƚ��>>���<�¾j>�i(>)�0�f���_=�3�=�ߐ>�Ö���=>m��-��7���鱀=����d���?G�!�ƿ��qa>.�>���\)�d���U�>hZ�<_%>	N�>1��>�L�T��=z�(�$K���$g��$W>C.�cu��:�n=��;�_�X�-�?R��=�I��隽����R��<�I<��?��+>;�+�<�S��E�<햳�|𦽊�D>�sP>��ܾ�Qؾ۔�ՠ���У�T��>����p�C����6������)>Lcj>��~����Y[Ǿ�6�>f�>a�?7r>�H�>����9��x��"�����k�0��3:�>R�(��+`��z�=g4���,�3�;I>��Q�ˣ\�%�(��G�=[S~���>�ƾ�?���l>^j�>ȝ�4��=E7�>�>��듾u�W��?���>S_G>���=C��������~���z���>Ea�=�R!���>��?��T���(>(��>!Eͽ$�>q&�>�$�>/��=-y�>S�=l� 9�̽po�=�$�=��?1�?#��<�H��� �*��l='�SUH���<��սJ��>�6Q��W!>�D�>3��>u�ὓZ>��"=F��pI��~�o=��>���=�`�=wK�;��l=g<����>Q� �Վ���}�I�;>�Ⴞ����@�(>܉>�1_�8�;����<���=���>I�4��?�)�Z���=�Ho����+��>sP\>�F�=����`䥾�=�	�>������O]�蹷���$�Q�d�9���=Ǯ�=���=��G�"z����>�;P�sh��LN�=->3�=��>> 2�<��4��>��c��sI����<���>�߾�Ѿ4�=��<���zֵ>)�_>���>T���A������þ�G+��M���I�mk�d��=E7�<��>w�h�RTH���G<\��=d)Z�����3@�<���輛�IN������A�=�M>z�J<�e��@�=�M�������l����*>Ţ�>:���G�6��>Hg�=Ġ�>n��>C�t��⽳Ő�
� r#�:|���|<aON�w%>��GwE>���Տ&��ݾr�?_">�8�<J<�́>�b���s)��������>�h=夲>�����.v��c$>9�A�?�Ӿ`v>�m<9����.�� 0�>{��=oK��Nʾ}z����?��eY��Z�V<�>�ǖ=;U�>\��>�<��`*J��;�:�b>U���ߩҽ�ij;o:C>uz>�>�Z	�KQ�>Ú�=�=>L�>�D���*=�0���k�o�L�k�=>�ݽv��SE>��">�8�G�.���=I�	>�>�3^>�M�>� �����0˾|^>|�׻kc�(1�>��=�eg�g��Xu��K[޾�n>� ?�<)�i����7�/=���=�N���>���>*3�>/Ʀ��9]�d���8�y\m�~����V�.;�=���>��Ͼ��4=y�>�̊>�������=!��>O�=�Y��@�=W��>��>�A����n2�a�����ʽ��:�����$4=)k?���=O��殾=�4��Ne���=�u�WL�=�A��!�=���>}H>K���Y���>���؆��X��E�A>/�=Qap>���=t�>�Ȩ>g����<�����>����Ň��>i>m:��[��,��h�>U��>��?��5>��j�g�L�?|�>�{�=?��>:�>�<�����oY��o���Ao�>��X>�-�>�G��|���V�Q>x�>)\$>�7e�׳Z��>z���kw�=�>� �>�yf��ݾ�O˾h��7���E��V�/>��ӼI��>���>����^����=\�S>
����	�>���=O�>zL�hX��S����>�z1�/Щ>�b�=V�>���#)>W������Ji>\�?�_>��>B�;���4=�O���h��ļ*Ɣ�+�>��|�7YI>�O�>ZB�>�L��)>������⽝��T\>���>���=M�n�E��=����н}H>`Z=_߽a�"=vd��h5��w��>�ͩ�� ���[��NCx����!S>�&�=u�>/�U�Z�>L��h����V���F>p���� =9%>��>�ɢ�})˾9U����=��=e=1��:�X�k���)�QkF>ů�>��<D2<���>�ࢾ��f�s��`7A>��>xڽ������=q���i�=~�9>�:>��P=��5��n��*1>>�u�����=�h3= "�<w��<�x�����ZG�=���>�~��픔�y�d>�9+>�Kg�[��>>���=O�����DO�=u���7'>��!�D4+=C=��:F>'{O��پi ��_�>��"���<��=�G�>���ӾP\���=��;�a�>dy��h�>�!��	U������g9>��彑�9<k�>孄>S�=��ۙ�k9��O�����>N>"?��~��	
�ϲ>��U཭K����!�>�ډ=��m>�qJ�к�>V�<>�DY=�N%�1L�ޙ�>�ST���c���vU>��¾�W��Pm_�j��>Dkh>�$ڽ���=��?Q�����>�Q>%I��^&>{A�<�=*�.��=��=����=
?�j�>� ;>��{=��޽�d�>�n�>O#�>S�¾��>>n�v=]�G���1����>A��=�5��E�= ��>j݃�0�̽�|���ވ>���=\�w���;TPw>1��P_þ8�{�F��>6�˽" ���EԽ�? ξ�~侶��ω{�P5|�
�޾E���J��=rv��W�>#W��I�:>av�=�*[>�|!����>	�>�$��r>Q�1��g/����>tQ�>b9Q��q���>�M���&ѽ�h��g����b>DM*�%�j=C�*��w�>����:$>x�����;&�>������=7劾u?T|�����,�6S���-B�����f>`��\��>'B<>;6?,'�>|r2?H	�=��p?��?i�F>[�K?!/�=?�?;�3 >��+���d?{﷼��>�>�>���q�>_,m<$#>8@H?�L>{	��||��?ɽ0A���i#�؅��=���m�>�H�>ԩȾ��>�9���G�>|�8<�B޾
HV>����B ��&�>�>i�g��G����R�=�T�0��=lcq�� �>��R�� �;YP�W�+?����qѽ�,�>�f?�h��?�?���8�8?DW�>���5�T>l�c>�����,k�*����7>�5>S�(�Ѣ~<}^�>��>� ���
=R��.w(���<�&�>{Y���y�>�Q0?�{>s�����5g�8�����ƾ�,�>�/�,'���fYB> � ��$=��
��>�?>�b���x=�D?[� ���>�u=1_�>/߾/%<���f& ?p��ڙ+��pv������>�A~��w2+���?.%�f����=n���>�&�>xm�#� >D��?�=��ݾ�+����>�T�{���㣾�
���}��mg��u]�<m�'=j��)���2�>���ߗּ��S�>��;��@}��F�>uE�	g�>:7�� �3�0{��ˬ=3懾ڿU���> 1�=��C>oӹ>�;��O�>&����u1��޾�w������3�x��=�c��>��>�i��#11<N���f��n��oF����= Q��QӼ,x�=L��>����s>�,����'??�?��a]�=FJ^�����K>	�of�>܇	>�&�Z�A= �w>'V
>�2�>zE�>��=ߪ�>wJ��ۇ�H��!��9<�!C��L:�>dp�>*�a>:L�>�+�>���>����3���Y?�h6�>-(5�()��
!>�	绑]>�@�Ӿ�+->\��>����*��O�����>J�� c���	�f�[=_�M>Rc�> �žJ/=%�>2**>K���+p|>f)��%]>&�f�V�����@���(�7�<pq>J ��!�}>��g>F����ӽ���>����> �E?�Pc?��>��=R�?:Ծ���>�wA:�c�>6�����>��?�*@>�Ϝ�t2@=MҢ�Mّ���Ž<u&>�w����J�R{�>����(�a}i�h�>TV��t�=��d���N>*X�>+��>���>Ǹ�={�"���?�h9>����X>6�-��[�>lݢ������>t�W>���j=��rA¼)���GDV�Dkj�y��=\��>4�2=��=��>�=(lʽ$mV�=T�>a�>7冾�����>��f��7
����I>(�W��ó���f>FQ?|�"�>�ľ��%=݅=?@C�����r�>��>��	?�*?�?T߽�����;��þۡ�=u��>���=��>ţA�Qh�>γ�>�K�����>w�N�*�a�}�J�^�d��̾R??�s�=cھGa<��?=���>�*��)�=^��>�>�I��_��>��M<��>}�%�@{���>z��K'>Q�?�����*?:G�>�K��	�g>�>>��>:�>Lؽ��?1qo�J@o<&S��p��X��>��=va>�e?�|�������?����+��:W?ro�>��N��Y��E�E?�!X=�~���O?����#�>w�B>ػ�=��>vǁ>�_����>�N7=��=�*�=��=��dN�on=|��>",��C�N.�iu���ݾ������ 4�����>�u�>���><�l��	6<��ܾ�m4���뽽?�~��󃇽�?����5ȾA�U	������f�l_>;�Ծ�r>���:��݄�U:>�|�ǆ�o��>V��>����Ѽ
Z�>h�=��w�:�B>�4_>ȣ?5" ?���+=A����=?�޾徳�����9�>ۭϽ��i>�b�=��>��{Yþ����3�'��
�>a�=-��O���7����v�Ӭm�;� �����E��6c�����S=�`�eZ�<��/�ֵ���ci=SR�#�|�ͪm�b*�>Ц�<	�콣�_�Pڈ>�����ྞ�r>o�5��B���_��>�X�O?��)���^��5�>�ӹ�;�M����=� s�O�ཱྀ������?�T�>� �S헽�=��H��y�<��������{i>2hӾk8���?�ߠ���}=�����0�=@PS�ԏn���.#�Em0>x3>P-q����>��ԽMK��wwn=��K����H�=w�Ⱦ�t��8�|>�D>D&?3�־��>��澳�>�u9<qV�^=�^�	>&ל>�o�Jf����=	��<꺖�񾉮�>K�>|S�8�5����t�#>
O�����őv<��K�M����=9s�>/�8>�\C?�>�x=RξV�þ�<���=���0Q3=��f��þ��v��∽B�߾��;��?��n�芾��ʧ����=�����T
�ѦԽ� >�^�=.P��e7�"m^�mX���9���(�������!�>Iy.>���=�>�u�=�[�>��\=�=w?���>\��2 �>�ڒ�Տ�=)��>�����̾�Y���]���=�􏽺	ٽ~�H=O/�<�˾-,?����&������>!�v�5�<��>>e�a?�|�;�R̽�k����>�
�=��}�����>��J>��>,��D��>���>,�$���<�.�=v�2>��p>����Id>|0�D�ٚ��!�>W�%?��?��?���>���U�V?���mH?@j?)���B�>��%n��"9'?�D>M^��[�-?"5��a#�C�p/�>Q�Le3��վ�'�� j=�Ɨ=)(U�xW�>��>?4�@��Ϩ��Rо]�g��?���l���㾤��=��j>�[�>��0>6n�>�ԝ<ܪ�>���$
��^�>߶?(K>K�N=���<�k�>��S>\�
?��4���#�Qp�>�G=���?���<D��=�BG?� �>G�B:B�?�h澑�W�i�ɽ�:���(�B/?Uˤ;�k�����>7��=Ρ>Y���(=>��>�i >�����?,�L=�����ٱO�>m�>q8ľ��ƾX ?��L>Z��?K�>�+4>���=�~���;g>�z�=��ѾV0�>��=�#"����,��>�H������&>��>���;�ɾ�->�`߼�ｾ��9>;T2?�8��L;,��>�> ���#��=��K�$",>�ɾ����݊>�:a��e��p�>Y�"��J����h�߾��
?*��E�=_�=<�D���#r
��P=}(1?Tľ.�O�o�>���~
�����D����x�>�ۅ>Y�<�a�>qV6?���>�侴CJ? '�>���=�૾_��=����$=��?�K>��N��Mƽ~y�>�&��������>l����. ����2@,��
������M$�=0?���>����}�>�>��G�s��[���Mњ>c�=z����>E�>Z��/�=�1�=�i:�Vx�B����=d���X�e�^���>AQ�wv)��N��҈>��=�=�+_�����c��=.�н?�Ͼ>k{�]�>on����a��q��T��<����ȍ����7��Kz�M�u=;�<>sy�;�S�?c��$O?M�g?���b�=����Ni�=4%�>�ӽ�7O���Y?0�N���ﾧ =��?���>�8s>��:>�I�>*m>of=�ӾQ�?[4�<�2��QyC�X�7<�E��ʙ�)\E��s>�J=~�J�D���ky�>x��g���vʾ]nJ���޾]��Y�T���&�%��=��߽��9j�p8M�ʤ���O��E?�&�	美�$?�V��S�=�h�=CAQ����2>;Ž�rh��=��>&�6>L�0�*��	l2�U�)?�T�V��3�T>�}�=N���\+��󾣐�g�P>�}?�P>g"Ѿ@�>k����D2R�C��>B�>�+̾�%\<���=k^���Wj���'�������,�(?=�J?k���v�>Mb?�BǼ����>/|?�R�0w�=u�O>�cK�7 �>��;ћ?#�3=&��=���<G�ở��>��H�Y�Ѳ�>��)=��=������	f�n���>��>��>�\�=���>?�о���'���г=~m��w��O8�>�]~>>8T��:�<L�N>��=0Tֽ~��>�� ?�3\��Pپqm���>�й�`��=.F>���>⿶��ӎ�����U�>��=��Q>��!?�t�>y�>����N>o�=$v�X~3=O��G��>���=»4������>���;�>0�`���7���S���=�7O>��c�iD�=o�L>f2>�Շ�e�վ�Z������v�E�C�#=MpD=��9��k����>B$>(P����"�ʷ�>2�ƽm� ��J���?C��>�Q�>�Ӆ>']�>��>F�=��^�A8�>��>{þC(ؾ���>��R�;5��Y��u|'?�G�<�>�,�=�p�=\&�>7���(�?�=��=�=�=� >���=���=����m���ͣ��ŗ���>sؾ8�Y>�G�>v*#<B�M��=?M����b���>vx�����5�o8�>|+���,�xTL�j!�`�>�vn-�_�O>$�<L>��>ijz�䈾�U?�5�>W���M���GҾ���������z>5�>:pt����;>�0˾��,���ȾݱE>��	���).�>1�<>Ձ���7�;��{>�1�>$�A=7�l>���>�5>{�J>�>��uV���1��H������>���>�eX�QN��>S�H>r�o>��>���։�=d�%�k��g=��^>� ���
�Ɂ�=�c�>�0�>Cۖ>�?N�>�yw>	Q��*վ#0>�Z0>>(����8�!:�>�:��b�=N��;H��U2��ޠ>:_�R�Ҿ�3����>��^?�1�Vv���B�>,u�>���=E�>W�@?~)=d���G��RF�=��>��W>�nɽ\�����=D�K�G�i�R�ƾ��N>�@�<U�_�`V>A�l>w躾�T�=[>(C�>W��ݖ?�T�=�X��Y�=g�N?�Q�=�����ݳ=>,>�2	>\%��uO>���������*���r�>�"ʾ�薾���>�]����Z�F#�>;���)���O��\�>�=G�?��S>F1�>�>�:>/������#t�;�y�=�ۮ>8�:=�+q=Xp
>pp�5�!�I�;����E�H>��K�}�)iQ�ʱo����=/(߽d}�>��k>	�d>�r��}P�>@(�>#�Ծ�����At�u�ž�� >�.�<�vJ>���=Z=�\:s��@����R�o_�=𜎾dо�9g>bʋ>1�?e[>	.?������Ӿ�f��"��@}���?4=�/??��b>SY뽷�>�.1?�wG=6�[��s�>�����i߽�쫾��a�:���G?,�����ֽL8D>0X�?8�̾<�=[��>�e�<��ڐ�<y+����W>��0���p�'����^L=�X4�g���1A�>���>��<��<��?���<�1�=�?��w=���>��>	�>.��>�i�>��=��U��tC�m4�fH�=$<>�w8��ka>L^&��$���!9�#�ѽ�W���|W���<��>�%���r><�;>ʭ?�����=��>���ZD����+>�P���ͼ�>��>L+�"��^��>��34+�e���~}>7 �|8׾�Xx>��>x����l>��%>�)���k-?�����þ�4>Hɤ>���=~$˾�t>2y>*�����}] ������n�!���n�xZS���޾X�e���½��E>ȰռܮF>�<c��w��>u����"y>�\>��t��Z�>[P��8߽��>]��h��a�'=��W?���LX&�'��x��>1�=�0��>���=ǌ�>#�w�}t�\�AH��/�z�_"W=��#=���l<>����<�>�S&��!���@">��_>��x��	���h���ܾ����>tj��v�=�>#���g�>�d̾�y+����>-d�>{�þ�K���s�<Ρ�>�g=��L>�[�>i3��i쬾���K1>�!U�Q~�<j�=o9ؾh�2��Q��#�\>K�>B����o���>/�W>��|��K��-?�@{������Y� ?�T��P"���	þ�7>B`�����O��uk<�Ɉ>�EV������ �>�C�=���=5̤�YK�T.��0����l4j>Y����(?}�r>]�B��ݘ�h����
�=�༛�b��XA�R�>z��=�&L>�����6?�?�>ZQ�>��=o^��
%>1_����:�r��LS�=VF	��	���k�>�2>��0���\�S@>ь�>��Z>��ͽ��T?����A�#�t�n2>�Y���I�b�=� �p���YK�('����q���a?}�k�5���W
�=� �>��N>��m��>��2�o�1��dξ� �C���8����ξ�5��V~=[Ij?$���A�]�"�>��(?�� �*f4>��2?9�=Q���RM�=�6��ZT�>o��>�Ʀ>�3��Oɾw]q��(� �)�˾_r�>qlM��:^��.Y>L�'��	�?a>�*(�p	>a�<�DU>ȏ�=D1���̾F��7=�2�=���m��'È>ꎔ=��>����)S?��_>�]e���=,����Q>u�f���.�z[�=�l>n!��mb�h��=/Զ>b��>��=�?��<�Jf���>g>��
<<L>�ͨ>݈ݽ��;�3��>ﹼ�]�=��?Zw���8��>4>#GM>4pP?�ڽ��4�� ��>4֌>]9������{-�=���=�]��0R��w���?��js<n�3��v��N�2�ܡ�>x>`?/#��(hB��>9��>��k]>L_>_!b>�%Ͼ�t��5/��Qx4?bm����>�-��Z�m��<�Kp���>1$x�4���o?̢>,R?��%K������<���0о�g���k�=�;�>}Y��X��=�=I>�=4?�j����*>��>�0�3���do>�� ��K-�����T������&=�u�����>|�v���p>���<��>kR?��þ%�@�7KT�ZP�����>��>G��=H�����>���8c�@�B����>/x���͋�=F��>ƹ�~BS�b��<�v^��P7���^��s������e�M>ҥ�&hl>���=�sO���?�]��lþ�-�>,a<>A���=I��K���C�;t��>o�?D)8=Vu+>�����>��?����w�r?�=���= w����[[T�yț�
�L?�����?�Hd�>�?������>?��߼L�׾7\m�e�o�դ2�b�>Y�b>!�f�����>�ֆ��b��s���>��/�T?���>o�>��x��Y�=��+�	��>���>I9>�ͩ��b@>�Pٽ����3<���>�Y�s��b>` �>쮾�y���x�X¡�7����>z?H�H=5$��Gv>�=�t��K�:�>Oc�>$X=m�~>����06?���>r(d>�	�<@�'��o�>�Q�;�W��=���>��o���񾈶�=�Қ>YL>f�>>��>Ƥ=`�>)�)?l��>�*�>!`
=3N>噽�s�=X]>�Ǿ��Z<6�?����"0�LY>'
A>�)�>U�>=���e>��>�B1��+�s��>݂�#k!�}}N��]�>�1�������p��
��>p�>�_��mI�(�L>��=�ڍ���^�Z2?Z%��/��o��J�>P̏�o�9�U���W���1e=o���D� �E��NA�>~�7=����t~>\��=_�>��?����=���>�,>#�;��<�G}� ��>��?�>�;/����>�~2?��
�hO��v>H �=W�'���S��r���>�.�>����p����<M��1ʾ߻=��I����=�<^��r��j�>a����i������|h>���
`�W6	?��
?tv�>�����)?)ȶ>���>��>�2?)��>�н�g?K�?�޾R����_>�7?,z8=�[�=�yq?�B>��U?��F?�z�;��=������Dx��5�=�Η�xz�>�!?1��B�9?�?�<lE@��:���)�>�܉����ڵ{�i�<�AD?�k��ߒ!��&���R��>�֎� 1�=ơ���0���?��{�>��9�uڽqP}=A��>��/��;?{9��펾wt�>_94?��=6P?�r>#`h�
�=��x?�G/������
>�?I�!?(r���&e�G�<�C���K��i ?�$a=?4>�'�>jQ"?%��;�0?�j>4>XT���8��p��j��>���oZ=���=�w���۹�J��>u
��h6E�R��;*�B�D�˾fB��!?�̚>�_?�.�>+�,�F�5?��Ծ [���>��l�>X����㫾�ؾ ����c��I�%���>Y�/?m4?���<+����Z���*L�>&�%�&�>�
>C��r�혡>�Ϻ����^��k��3/����;��o�>d����ÿU"�3=>Qͧ�>ڛ�Tܯ�^{���6�l�����=�i?���徉G�>4t����?������>�:�o
?�D��FF�>���E�=;H�[�F���Ή�3>ö#�� >�
�Gm_�M�s?�<ѣ(�>
�����>�t��z+{=ʽ�|��<���>|�=o]��{�>6��>�SY>P�>ہ*?1����%.�i��=��R?�>Zҽ�鄾�9���>}$����.��E�%�=02�<|C���]>��]��ڬ���$�
��>o���u�۾F��D�?N�?}�k?��l��>�?}s?�^G��,e�ϋ�����E��%�6;�8w>u�==�.=��H?'FB���R�IӞ�V�����>;TX?,�=�������>�ͳ>���>é�=�2?s�>.���UV��Ad���>��=1������l=�	�z��;HW>��l�S�?�߭��W��0SȽ�`J>��b���>	��>�W	?���>��E
?�A|��v�=�h>�8:?�,��$V?���>�>Uu���g>9�{��fi>I�.��=!�JO?��}�>3.3>���Iv�O�?�9
��cb��P��z?���>�d+>�q�����<b�w�Ġ�����=i��.y|�UW�>�Ak?��ԾD4�>?A�s>���&�>��q�bl�>X���_
}�hþ���?�L?�M-=<�=��t>+!��>2i��IoW��}7���l���j��>�J�d��<���=��4��{��]C��P�G�_W����>�M����ξ��A��Q�?�4?�6�?i�<�	�>�ᖾ�;��r��p����4?��?Q��m�5��W�<O'��c�>��f?��=Z��>
�Q?
�^?��(���U?��?D�>;�;�$�>��=A �>��>��ȼ�/�~[�>K�~�X��>?�k=��7�C���.ԍ�?�}���?��?�L9�&f
��,�>���>GV>��%?��ý�l�>#;"?��?���>*X���'>���=u�Q=6Ʈ; ?��=>�;?�R�>b�R>�� >������=�>K��9��%�<?AҺ?3�N�ڧ>�[�>G:?(o�>�>1R����>�#(?g���t�:?x�Q?E.����J>��v�/��z'�>�8v=KQ���&���ʻ
~�k��>J��>�0�>���)I�v?W~#�iX�\R�>�B̾�t1>�k�=uȋ>[��E?�I>��=�x�K�f����=���;YDľJ��jM���l��R�>m��=c�;=s���>�4�>>��>���,U��OV\>�(L?�G�>H>S�>KXE>�39?�~���0���>��B>�]ҾT����I޾v��>�nٽ8����ھ���>#g�fžԒ>���'��(?]��=�y��x���j>Ds6>�C�����H�=O[�>��'?��8�ik��-*b���>y/�ж�|˺>�(=��~����>���=S&s��
�P4d�(��>./@?�>u辷�>�h?��l�����;���f��<ނ�>˓6�����L؛��a��򢽼�پ��E���>i�����辏�B>�� ?�$���� ��S���>K�D��]";�1;?چ	>}�����R����u���h�0hZ�0���&s,>Ϣ5�M�׾Y��m�վ1>�X�$��f'>�c
�Yƾg�>�Gp>E�
>i8U?�X�d�1�Aց�TcD?P�U��,<���g�/�>��4���>s��� �q>!l?螧=b�b���?����H���>�}O>�S��΋�=������$?�񔾐�c���>|a?0�=��>��|?� ��\���<�>� D?8"�Ք=k�=���=#(��X��c���В;��l�cWm��!u>���=�$=za��D�#?���I�-?�\>�9�=�C��+h�d�ľ#�X�2�¾�G�te??���?%B^>�5��q�>Eh�>ț�>�y�<?9=\�>V�>fu��)�3?[CH?�s�xN���r�>�Q����X�ξ�qľ���S(?�kX��G�R#�nt ?���=�(>���ҵ� ��=g��<��F���(?�뢽,ב���a��BU>��;�����0�Y�/?j>�7$?|�{�>��c>�h>�o
�ͻ�<�q�>�Ƅ�#�<�s�>�k��#���t>{�?�o*?�w�>���׾�>z�>�~�=7[L?���>�|��ݻ=�E?|轍��>d?�>�h���Ͼ
�|?`4>s[�<�3��Q޽�j�ܮ>߂Ӿ�ɨ>V�
�T�2>~���Zv(?����v��=�y���l��>fV�$�,�rs�|�A?	�?���>2�}�HV����T>j\�>�t5�	}��ۚJ�Yf>��8��?�\����1�:ٗ�Q�޽,��:�>(�f����,�?�G?܁�>�*0?ё>/σ���">F�<�D����1��ӝ��0? +i?�z�u�`=Ғ�>��>y�>C�ľa]����>��7?W�+��Z?odY?\G��&��=����؈�>}�	��V>�ǀc>^�?�'�s�k>��?R?9%��8պx��e�>R�<�,�>o��房dD�>Q������_���5�&����>����4���A�>$����+��5�>z�����)�Y�۽a�ќ>υ�>�I�?��� >��B>N�>=wJP�X6d�(9>c
*?��?��>�h��>*\h���=�?�@?�A����}�>�?ǽ�	?Q�Ծ�"�>���⟋��^�mk�>�SO>n��l�>�	�>���>�u=[҆?��>�������j�'��`<�"?
�*���"�K���ͺ=_���6E����	���e��l@>�d+>ڷ����?��ػ>%{R��a��V�>�/?��󾑬����>|Rվ��3�"�-�q����]<F>��V�D�"�z>p����M�M�]>���=���>Ծ���>���I�5�e%(�u¾>C��� ���=�t�>��>d��=����H	�Y4?�e��c�b�п��|A>�Y��7{V���;7��!����F��; ?Qy�=={=��	�tK�>� �>?�=�A2>��?�=�s>��?�]�>1*?�
?��T=YE���"?6�񾐩���\���a_����P�=�̅>�0�>:i�����=�d�[Sq?�?N����jF��ݽny���[�H�}>"c?w���⿮G�u	�>x���Z�߾r����g�ÆͼZ�{�l
�G�?w`ؾ�#�Nl=Nx��:?���I���{��t2>�t?�ɾ�X�o�?���>/�񾡣��`�=�ǌ�>�_k?�>K�<���?��1?ط>�[���=��"?FѾd���������=�o���.�������=��a�>J��>��?
>���I&>���=_s>z������>4�!��K���ۂ�I�K��Hν���=>��Sz=ǡ=_t�=�E?�e"<�6���>�?9ݹ>���=���>>}?�8�>��V?�Cf?��'?���H%�>�׸>q|�>.�f��>�9a?}o1?Uv�>-����>ָ�N{v�����������v�=1)�>���>��6?{ �s({=jPc=��g=���>ϋ�}K@��7��ך�=`�ﾥ�=����%��>�t�9�V>�Z?��L�U��=5�&?lZW?v��>c�N�h� �����I��|����A����>3 ���>�<	?�%e?�����R�=H��>&��?%�\>����.��n-?#�(>k���=p��0l�<��[�覢>���>X��������>EN�?ఢ>� R���:=j���9�F>���]$��
վ�@A������U��lG����2y�>7.ӽ�W��$��>8>	�?�V �d<;�KU#?���=���?�x�G�X? �X��#�����A?)�����F��@�#ʳ>�&�>95�?�8��#?�����x�>F񙾋1���|�>�ϩ�%A��R=��>�ӱ��ɯ��=����L���=�����hha=�_ʾ�v���'���^�<�K���3�ڞ�>U일R��q@���#?_(��m����D��/?��-?ٛ�=]���"�=A#���X�>9_>]�Ě>�'?�	�?$������o?DCG>F����¾��&������z����?�5??�)�(�>*�\�x凾םu>Y�M>Y�`��3�$�^_�>F�����=l��=+i��AG?㽳=]?��>yU>���������>���C,e�p�l>)�>��(>��P�5=�JS�!i�>��>�C�>���>إ��;p;��Ɗ�;�J>7�T=[�_����>٭X?�9N=�
?2a���g?�=?�:�(��ҽR=��-=��F>1�E�8�;`O��f;����Vg*�'�'��=v�\���;�F��>H�>>�>�ĊA��v�>/ˈ?�]׾`֔��e�=��?tm�������0�^7?+��>YTp>�(���[m�s�����<<�>�a�|���ϐ�
|꾕�ܾ��&����B��Ɵ?��������F=Y,����>	��>(n�<�z�b��>f9?�8?�+��\�L=i#y>�L�<s�?��_�>��}�]0;>G>c��>��~����=Xړ>Ͳ���Ǿ���׹J?�,?aV��TF?�M?",���&��Қ�m���A���D��Z��?8��Y.�;����y�p?�
>V	�S���/�>k�D>� �d0N��½fiq�/�>��f?5d?��<��!��u4j?�>��s߾Qa���m��ꎾ>{1���2��^�=v��?V>Q<�D��R�羿�>�����1����U��>Gk�>m�?��A?(r�!(�����Hj��� ��
�� �>�)A?����Ѝu?)/\?��>Z��= ��>aa�?��5?�)��D��Y�>�ԥ>|��<Rf�=��>�5?���:�����>|K�?�#$�L6>eG>�(?�60>�i��Zj��S��Rv?�M��!�Ͻ�S?T�<?��>�^h>{����>ŃO>�΃?-�>65?s�=D�?�L�=m��=q�>3�R>��>�q\>l�}>�) �ݣ�<-ؽcF1�`�R>�2��@:���	�
vJ��Z>Q,ϾTy�>z��>�x�=7q�jσ>l�>��?H����>N?D>i�X>�t�#(F>e�?����˅���־,��P�`=�ߐ>�_�<��K�����m��gh�����>E��>QBm>��>�c�=�'��lQ��?��?҇�?,>M��?4�r>�H�K�C�Sen�����b�l�+���W�Ũ
�C,�n��>7+����>�k䄿��v��/[?�?*`=7ڷ��cK?v�?���>D�_��"$��O>9G'>_�������������>є�4��J>˺?�^�������)��?�}�G�a��b��۸�}J��Z�
��7N>e��1'�>��>��
���羇6����q?��@���鼐��gz���X|� �=Qv=���"c�ۈ����E?`1�>���Dkɾ?��>�L���:>��p�����x��>�ȡ�%,>V����>_����D�p�(>�X���_>��<��Ѿ���4���E�=�y�=�_��/�x��?Zd����B��������>���>0��=.��D{p?uV>D��<K���r�=^^>;����Ύ����E�=T��>]� > ����#sE��@���m��L��k���2���>[c�>#�D?�`?�M���ö=#�%���A?X�e���-�{ڋ�<*��5E>W���>9�oܔ>l=��_?���?����E*��5F�dW>)��>Bi>ע6�.�g�+����=s�(�>h��C�>���>Hj�>��(>C?	7���v=Z÷�Aɦ>�B=�Ry�U��<��=������f�ʕ̿�4�>q�?�k0?���>V>^_f>z�B?ܐD�A��>@c?�����l��/�ݾ�y�� ��i���X
����پZ�I>�?��߬���>��I?��:3�=���>|(�?Cf�ZK�=�m>;/r?�5�h�>H�>=���=*W,�o��>��><�E{���<<����C0���ܾ�C����[��k��=6(�>B��>T�v?�7�P�ھҕ����>��0���t�?�O�=�����YR5?�u�>	ƾ���8�C�_���<Yi�<¯�<x�����	��"ؾ&�� ׽۞j?�!=�_'?��0?�S>T1O���>�i�?@��>��>�#%���>�H�;'��<��F?{�f>��?�U>�*��fM�AK�>y�k?��?�{���E>�d>�愺R����8�>��=4k&>�¾�Ӿ,T�+�p�̙�����>֡�=lG>�'?�<���=�t>?�8|?�>�Z��[��ظ�?��AC}���� c�> D���˯�d�����>p� <A��>vT�>G�>AD�>�J;�"�>�ID��>!.̽���3z��y���ۺ���='=���*�>�i#?��=�q��O�>K��>boL?�.>%Q	?bj�>�h>Li������[�a�%�j=�=|*�>�	>�t�\5 >��
�32?1�CP���7>�!?���pD�H�~>�:?�!�>VA{>'1��s����$U>��/���3�^����w>xc+�@� ���������>gX����o�#���
Ӿ	�>��������>���u�=*��)�>Oѽ<ɭ>虖>4۬=�vc��]�6#>>���>�J,��[���w>, ;?i?���sy���L?YD�>����.A���\����>f�<>��m�W/���?}V?7
��g�T> �?��n�A�W>J�ͽ��?Z@�<���;���>�]��xs>ee��P(
��#$��$�>P����DӾ�����=����j���ؾ ���۱�>brB?�(�>�x�>�q���\����<���>G����#��#L��G
?1�c�}G���6�J���j����>G?y�������=���>����X�"�ԧC���>�����,���?8�>Yo-?A�:>���E{�>����/�r� �1�>_J+>C#��v��Q.���=t(>;�]��{�>2�l>?I?��m?<�E?�y!?�O>ID�=���=9T�<�%7=?�ѻ)�>_�o�h�Ǿ�]�>�ZE?D�Y>\���%��>G�>m�t�����h�f?x@y>�
��ԕ��+>�˽V�����os��m7>�	t�%|5��&�>,D�+~ �.�#� i[?�9z��+��*��p�=�ɑ��L���
���8��
�<� �>���m��9Cu���=��"���>AA?�>����5���.�C0?x��?�h�=���>�ۨ>`+�<�j�?b o>��1>�1�=ه�>/��fc��k]>�Z?�U���y��_肿e�>�L*?Ot�=z74��f�=�;�>���ɽ��moI���Y��� ��nH�&]��"+?�{��!>tYB>;R?f�>�D�>�O��$�>t޽_=+?�dX?�>!˞>>�V>�����>���@?�>��?��?���>*���J ھ�l��z�-?/�?��>��K�^���ܾn+=����C>�oľ����+�>�p?����D
�=�w?z\�������ƾ��>G]'����|�$���V?ې���Xz�^?��W���=}�Ｔ���N "�M��>�Y
?+��>K����ؾX��F���t�>3n�>��?|�C�p�>PI?��=��>A�>)�m��3G>\���qu>�۾ȇ<:�Z>*�?�@�h�:��>�>v�a>���=ju_��'�=X�1?��o?aq[>�AM��v���Y���Ƹ����RW:>O���#��Sɾc�� ���.!�=޿T?M���(��;����>$�!>��>/ ��5�>��>U=�>�r*?��k?�Ʌ���-�)?݉�?��=��I�X̿~1?�H���<x;�9=`n�I�9=�h�aq�����L���r>�2���y��;�Y����-\��Z_>����`�;�Ž:�|�7��>�z�;ʞ��A��O��t(>�6��ҁ>*���$׾�B�x?�}g��'_������>�F�  �>`\>�c���>���bqO�B�þt��>-$'?�d>ۧ�<�l���R��]Lo���>�
��Iz<�8����1>n�̽����yT=��=<W;�G�D�F����>4���f㪾T�=zq�?���=MP�>�e??0�>�$�>�X�>�&�>j�u��� �j��<6����>蔾I	`;-u[>� =L����Ծ���>��=+c
������z2?O�k�'@�LT���*��˧;��<�z�>��J>+X@?g�>h�G=�c>+N
>";�~	~��2���g.?��>�l˽~_c���;Q�OS������A�=J�
�H�9��s������%.>���>�þ���x ���a=?T�`?��%����>�2=�{���s����=r݇>4��K_j�
���繾§�I�m��=UѠ>]vR?:��W����j���Ͻ)>�9ǖ>��=?�Fǽz�?m��c/�>>����=����A.�%��<�B�>�4�>հ�<��x�����ӽOe�>]S����t��BV>C��=�]A?���;*�>fH����ݽP��5ѽ7v��f�>�2?�.�����(�*>��f>�{�>��>A�l�-�ǽ{b0>�&�>�+O�M�5>��?*�=��۾D�\���N���˥��A��9S>C��������=:g>�1�>&�>��W��L�����=֟>��Ǿ����:>��>��=�=�*Z���T?7�ʾ`���վLw=��9����?[~>6�?1!?���>O��>$l��K����F���M��U�>7^�;�
>i�	��
$?�6?�K��LB<�:�>k�>,�c<^���kg�?�W�?U:>���� ?��,?1��>o�ھB+>·��}݉>�$���#�h�H���|�e���<ھ����MӾo�8?�Wc�s�n�Դ.?�^?ih?��b>��߾�_y�ps�>7�^?n��=��>p>��>{�*e\>�J)>+��>�,&?�#q=�"���-�h����P���(?�>�Pi����*?ǷJ?+7�=�*��z�,?t}�>��K�6�x���>ʁH?
b?ھخ=�P־�/ܾ�W�=AxϾ��,���;�s��e���辎ź=���>򣳾��LX��s�?qR>k�?�?��?~&���gʾ̔c��1�>
a�>[Q>��t�C�P���-���#�����&:_='�j>�Mq�ov��n��۽��t������.�gQܽ��Ͻ1���H6?g�>6uH��'��W?�ᢽf�ﾬ��=�?8��>{O�>,	#��*$��荿& ==�T�\��/.L>r�?)���x`]��iG>���>8A�=9۾����3پgN>���=��!<��>�#��>�p�>�b��2��9>k�}?��=}���P�i���Y����*��1˾�$�=\>)��c)>+����T�>��Q=�t��`lL�|�>��?X�߾���>��=bk/�1_??Vc���>��>�X)�����8���$�Q�s>U?<Κ���\�~����V?��������ܻ>�Ѡ>��k>�	�$�@�wX�>�)w��g-�1s�>��>�X�����:��>6���6�%�˚�۾���>��R>��
?�^��o3�i�}�J��w��d�=/�>��*�&Z��ӆ>H�^>�j> f�>٤j�S)���ξ�>���>B����>��@?��̽�슾��?Պ�>�X_>�c�=\��& ��MM>��žձ�6vv���>J�9( ��t��{?7*۾�D?�U'?y3����a?(�?/ʰ����rs>t��> DL=�W������1�/�`�>
�������:�@����G�?l�>�F,�1i���>yY�>|�[�ŐQ>M\��1Ռ�#Q���F���q�+Hp=hE�tŌ�^(��]#?��?P�!?�<n����=n�F?��>	�7��,>|�?��,=˖��-�>IF��JX�L����׾~Z��WQ��
c>��	?�&e>�s	���K���)������</1һ\�? �Q��p����<�=�N]��ܭ>�P��|�-����<�T�>Rt����=�	�>�W?���8id��Ā>PCڽ�e������/?$/�=w������������>F����a=�et>Z��?x�h��=���>i��>��='�=�\?B��2��Nн�/@>?!=`��P?i0�>�*�ά�b=�=nc>�.?���>#����TU��N�=��(?��>U�3�9�i���޾����ddO�-�ɼ���_�O���y��>7�H>�h`==<�?�>�P?`��>EMǾq���3��p穽���>�->yS�>L�=��׽D��>\e��,R��m?�Q�?
�?җ�=4�ƾW�ν$��It�f��R��]F������c���>��2?��>�`��R?���>��r�dU	��U�>�v%?�S?|=ľc]F>û���ᾭ0���C�>l1�>�ڤ�Rw>߱�=��=%�>)l�<n](?�x������Tq��]���>�����Bx�>�d� C���a>�'������X=։8?6�����i��Y��>�ץ�9�>���>�5��{������Ƞ�_�C�kb	>��9�V>�Lw�K�>�j߽6���Z���g>�G�>�ѹ���ʽ���=L��>�a�>>�=R�ͽ�L���6�'�>�ۍ?BԆ>����A��[�����5g�t���>�߹>T��J/�<��et6?��X?� A�vd�>�(�=�
U���e>~7>���N's��)�>Ja8���E��[��@�<�i,�W�þ��2>�W`?a�˾_8T�ts�t޹>Zh�����>�\�>��>�/�گE�LE6����>B9��ƚ�^�����<?>��cHx�?v۾i�>ᶹ�䤣>AI�>��W��tp�[v8��M?�<V>���b�L�d���)�{��(
>���=�?�Ej�>����y��!���>������x�)>|��=�`��h���c���?���YR=��C���>nk>C�>�F?	�m?IE-?_
�>�r?%Eu>�h��G�=?���A�>5v�����~*�M��=��Ͼz��� �=Ԧ�?E��>=Q3�-eR���>8�a=P�����%���?Ӎ־I瓾Z�&�X��W0��E4/<��>�2�����n��9(�~�Z?Y19�,&�������>g2��Pbu�Jr���x ?�O�;%zb>p�:>H�V���y���x��N�tde>Q�)�?���ά=y�<
�3?뿞=��/�|!Ž�Z?��W?Yu�jg�>��>!�2���?���^a>��;�B�ɼ	�K'�����b�1�J�[=<G�oM�=��>�Z ?�l㾚���Y'"���>����ۦ#��\>O��>A[#��ͽl�$>We$���-�B�0N�>#_5��l~��{(��M|>�� ?�l�>�ă=��>��a>Y��>65����>�?j�>Ζ��3�?N��>�f?������'H�5*>�&�>��=\[��5>��g>_U8���7�y�������I��7?�a	�1�L>S��=蹅>94���� `�>��=�1<����С?��$���>�]��F�>�X����=���=wH�>-Խ�~�>(s>A,6��
�p�>�9�ǲ�=��wO=j�!���콬"*?�s=�~>�?��=AQ������PI4?�ڭ=f+ν"3žnV,?�rv�ix<ڙ�����?YU��&�?U�= H�����=�1?�t2?�S>P�=T6>\�>&�̽�����D��:�>�n�2y߾�w%�VU���k��C��>7��N�7�����#�Q?-X���@=�G�=M%�>��>>���9u ?�m3?��)>��=nZP>�ΐ�7�?�p������7�?uн�B�ݾ`��>�>�>H��>P�>�\������?b�	�٣��T'�=��/��==>l@����U�H.?(��=E΢�
�ڽ�	��̈<?�H����X[�R��_�����\�P���Lj>/G�>����!�<�B��a�f>^�a<;E����>��o�f��>�=ܾ�)S>�x�=���=r?��>�����>�o����?KO�����no>�N7�5�>Q�.��ӆ<�p�=�U�>���(8�$M�>s��>?�������V�>#�>\L>u5M�F,�>�l=?���>{Uf>�Z�>�ľ~�+��"�z[5=������ܕ�0��>b@��u���F���z_>ɾ�>���}>��.=/J=}W���<���� >B�߽��ݾq�>M�#>�i�>N�
����>�ۖ>��=X��>���_���9?�Z�=Zn>1Ğ>�搾	�>rڢ�s�>���=�7>Dna���u�go�>E�>���ቪ���>?0V?��>��7��'�>%m�>�M̽q������3>�3M>'~c����m��	F:��Z�;�=�S�>t�������i=A�W��ך��a���簾x�>I���#��>l�������6�����q��>2� �>�����>K^�>k��n->Ru��(?4?e�AE�>�z=�p@>��?O/���]	>i�˾��	>:`�>�H+�Z��="�>���o?�o1�'��?���a�?�,�vž["����>�g_=���=��8���>P�-?{���8��=�;M=@?ċ߾�����>�i��m�.=��p�Z-�>%?
mA���`�X>�U�>l
*�TW������˦�>:�=���B>X��pB=[�N>�=��
��xd���Ѿ,���d��T���?M>�+�>��6���>�@��颾;���Ւ�h�>`�>��>4wr<5�?���>�QU>Qã=T/�>4�6>-�&��v�>G����5?:�,?���>�(��1�>}$�>��C�]�:�7p+<?�X��x��徜Կ������GR�7��8��̶߾�B�J��>Z�?;e�>��=�<l��>�4>w`���)?�y���Խq9!?%�4>?��>N�e<�Ì<��>k�D����>�^�=�����>W���ȿ>�����V�>5ď��z��w�?:��>B;�>���(Qa?�.�> u���_�l�> ͝>�K7�����>�^?*	G��=��Ӿ�bٽ:�F�=��i��Z���pB>��=@��yY��xI>O�3>�.�<	e�����>O���=C]�<���7�/��=��^>�y��̄>�n[�mE!?.Fr��I����;j\	?��C��y�tz��qнT�T�����?1�I>��'�ipM>M=QI?1@�]��=y4�;Cr??�4�R�=|��<��>o�?�������e�?k
���=AD�����>�;���u>�냿�Q??)HӾ������`��j׾j��=_N=>�>�-��þ>pQ��t�>&�.��g> ��=?�&?[�/�.w)�V�=�����Y۾<����>ҖW>F;�nf�<g>D�?P���{�����We?�����Sy?t[�>U�_=&��>/8	���"�C��P��[4� ���Ѿ�"	?gu��$]z>�ʏ>���b?'�;��R�	�<��>�C&�z�� w��{?1��������]>x$�>-�)>c����3q�����<���+��<�ȟ�u�:7#?M�>�a�>ʒ�<���=v�>��Sy���t��I��>��뾬�>j��EI>�R?���=-�#�m�t�q}�<g����.ʼ,�h�^�>9{�s�4��+�OI?|�?��>�Hs��K��Wa>�1C��%�fc�>�?P>�CʾB�����>��=q_<�x:��g�>&��>}]?>�Y>ip>��0����>�w�>��>�x���4>������ӾB5�Y�Ҿ�h->*m���)>�^>�<��e���h_>�Ӽ(�=:����$�:���ܫ+>OA����=���1V>k"��X�9>?*�'?��"?�7�s�?G��>(]}=�۾�(4>�E7�*��=��.��=�X2=]��=�v�=P|���N>�� �i�� ]>Y�>�%�=�9�>��Ⱦ<�	>s<;=�o�*���&_>U1B�?��>Y	���>�,�>���%-Ҿկ��+�&�.`�<-@��|�o�>lo<��?=]�=��bB?�R�>i���'�.�agu<).����\ �P0�<�"�>{ʾ�+ν�	?�P�<"}?�����vi??Oq/?��>��?h< y�������fŽw.%�[(�=(/����>Q�]=w��=��=�W�>˃���{O>)ݗ��nK�cg�>C}x��9�>���C�)>$ƽ=U]��!����� �܂=&�-?�ɿ�t��b��>��?iΗ>^)w��?��s>�[=�z<��>�tվ6)�>*J޾��&=FG��rP�>�_;�>w��>;�F�	��&?��
?h\`=56�>ޏ���>����<�b�	>��>OVA���Ǽ@?��>��>��[�E�X?q9�>��!�ӆ���m�>a��>�����E�P�>��?	9��m��ߠ>5	�5W��pC��%��>U(+?���>�엾j��>��?%��$Y|=�-��)>J?(���;�>�C;��Y�����F>~.B��3;��>؁�>b(��Đ�����z�=O���Ң�C%�=R���P���Q����
��k��>��>�p��� Ͼ���>V�4?kmb�[x�=_Z�I`&?SA-�I먼B�Z>eL��{)��u�u=�Q�>�WW>�,;��۽���=:qC?>�(#�>g[h�mT?3����3���=��I=t|��w'��ωe?�=�>b�#��[�=gX�>��n�����ˏ�Bۈ����'�=�w��t��:׾�W>��m�����ǯa>u�>��w�μ�/��<��(>���d��]t(>�>�E��?��A�Ծ4]�>W��.���D�0>{��>Z��:
y��a�=�p,>��Y�B�
�.�J>,�e>S����>��z>5Ǿ*�?��ɾ��>�<x>�E��Z�>_��=�~�,��>\�|�dŻ?y�>*9S�����E�ÿm>7\����<F�>m���������=�px>���	�ǽ� �>Ԭ�>���>^�>ɷm>.!�=�띾�)����<�P�=�̓>�>(>č�=��D�$��>70>�Ӿ�Y��0�X�?�ӽֶ&��oýAH�> ^����>[i��,��>S������=ϋd�	D�>xi��zT���>@��m�>�A�=R�q;=�+?iɾ+�>}�p�)�>���>c,0�
�3��Q��i�L�ȸ��pu>-�7���>�L�����=R�>A\]=�ɼmM�>�缃�%?K�V>.��=��������?k\,�lnA>���qۆ>p�B�	ϫ�qn�=�6)�3����p>۰��t�?kܒ?�_�>;��T�=*��g��>��#RY?3�c�JR���������((�l�辙�R>uU.�r��1�>��p?
�=ڰm?��8?�qA?,��>*��?���?�v�>��v=RG��!8�J��y?ḁ�	�?G���P��׎>���,�>�DX�4�?�O>/��>o9]���Ҿ�)G�J%D�����=F�>�`?O�@?O�!����7K>=��N8?����w��g���I������ླX�>EN�?a���c?��s?�ғ>�r���>�= �>��(�*�ʿ�K2��pp>�(;��>��l?!?��?ԩ?vC�?��>�<�<]����4>��>�k���?���l���7?p}2? Λ��<���e�?wkl��r�=K��<�j��E�=���>��ѾO?�A�>��O��s��:�>6���]k�����O4>��J?��k�t61����U��?�dr>(����!���Ő?uݾ_�r���ɾ��D�*@Խ��>7�>�g�>(;+�wX۾�c>E�<?X-��:�ϗ���??P_>f���hfR�\x>{��"��ݿ�ѱ�������X��3�r�$�M�S���36�`̾:��>i ?��O>����հ>��?,%�,�?���Me;��~�=��P?�o�>% ��|�>��T��H>���1��C�?�N?gQ�=��@����gӻ>?����*H�T6���Ҿ %�>ORA?+�=���U�?(�L����d?�?Y������>L;F��>X������U��=�&���a
����ƾ|p��#�	Z�<�$��$�?N\�>D�>�i�̗�?{�>%���ܾ��?C�������>�u?�8?�t����=��?��>Ç=�5���?���Q�:��C�>"���9���7�>���`�a&'?d?���:I�9�l?�D�>݄���/޾O��ωr�c�F?􇫽rK���H>���&Z��v�۾֯ؿI)ܿR��mo�깮��32�y�+?f"ؾ���0�?}���K�_�@?K��>rV	?k���}<�À3>ps?�*���v1=�%�ɓ=�6����C�h��� ?��.�Q�%�R�ec�>��?�J?�2?P�?Z^�><��>~�/?��I�۷}>ڒ�>��཈RO��_�?���?=b������<�>V�޾ (��*�a�WT�u�_�	�G?M��>�﫿�O�'�?�L���O'>ec=<��N�~�H?!nH?U�:����;U�#?=3W�E4�I���&5^?��>Z٨���ھ�	?��?����F�ﾏc��^c��k��9�����{f?���>�� ���?4�?�1��24����>y�|?�m?U��=-���W&I>o.�?������_?�M=�N^�3/"?g��>ڌ�2��>�Ϋ�c����*��x���ھ�bx>Yp�?��>��%>n��>d,�n��<|�����>W�>�I>p~��؟?h��>��� G!?3�>J����G?ML2?X����Q{>W�>���ڕ���E�s?�Z߽�䰂;��g�{��?���>F��?! ��d|�?dL�f����ѺC�8�0?�hD�u�?)�M?w,�?�#@�?p��ٕ� ��?ִ$�y�7?4��>ؘC?%�>�[���-��D,H�t��=�<?0��>� .���]7"?��w�h/�=��>�=�tO{�z?ݒ?m奄ր�����? ��>��Q?����cEʾ���{ �?��(>r.?���=ޏ?@˾�_��c��i�=��=�>��$�=ts���C���
�l/~>����qy���ཕ�>x��=-mC>� �>@��)lK�+g%�2�&=��쾜E�>���V�\�>(ɪ��i��Vk��X>�$�#�E��zO�(aH�#8,���?N��=�s2?̨j���=^��?á�?�Sa���Q�.S\?k57?]�t�Z����r����E>ߞL?5f����t���h�>�@���{�*N���=�n�?4ٓ>y�b>���?U=�.�=��~	�>W��<�\?ϧB�!�����?��?��Y=L����Q���$r&���T������y��ޓ�U�����	�.�?l=��O�>��?Q�?�w��B���?r�f?dK���ư>�=<�%�_��>y
/�����F{��;�A\w?}BC��l��o%?�U�r�Ŀ�m5�:�'�5��>��̽�#7���=^�e>m�&?�;h�Þ�>p�p�!5)�>G.�����h�?C歿>rj�Ɛ���i>�	�����-����+�յF���;Q�˾�F�~N��<��2��MȽ86�?3��2�7��>96?�\f?u�A? =�����z?_���??p�y>G��q����=?�kN�ѯ���!@��v>�G��Gz>B>�=���<��a�
�J�=kԾ��O��:��QO_��[X��l�b���� �uň>f͉?W��� �?�"�>z��]�O�F�?�� ?�K�?8'������,U?<O�?���>����&>�z�*��>X�=x;
��E־fm�>Ǫ >��f>�y0�)@�>/G���Q��_��=��R���9�����wdQ>��?qrp?��"?O���5$��s�?�Y�>�^�(I��@?5 �?EN���$?
��>�q�?LI�>�$c�^��=e[��w��ۍ�ͅ�>Ǆ>p���k׿�
)>$�6���>{�޽���SB�>(��7��<���H~?P؁���V�Ǿ=\�=����]�}��-վ;z?+%>�s��!�t�4��#|>z�3��0=�6�=y����R?�˹�
a?�]k�g�{��6���T?��??��>s�l?���?�x�<���=�j�>�t?�p?5�Z=����F;�42#?ε?����7A?q���kl>-a��'���	?�9�>��>C5$��??��z�����4E�!�x?܎=Ι;���&>�������0�w�c���_�~�?F;?�A?�1)���˾��?��h��KC=I� ����>�c�>��='L?H(?�rj?�<�?���1@>�fǽݹ�=�	�3/���J?��d>S�	��[�*�?T2��YI�"8����w�|�G��{*?u#?�m>�N���m?ݟ��.��>�6�������A?#�?��*?�|��}�>=��>A�>���>�\����?& ?=�$�hJ�?�&?>�?Z�0�O����c��n�?��[?k?y	�>�Z��41��`˾�#?#R���Jx�sL>���>[�r�<U��,�X���(��>��}�V�&4m�Kl��?�z��]���U�?e�k��>?w�?��=C��&0�Z�e>2+H?k�X�w>9�T>F��7�R�?g��=B��=�򾁋�>TԌ?kЉ>�(���?���?[~l>5�M�AH��s��+�?�Tǽ�b�kNB?���?��D�c���l��gt�?HO�>+�4/��"+�=���?�?�4V��?J��xK��!#?ç��BP���"��=�u޺>��a>��+�����pS���=������>,�M��-̾�u���5>?9ྷ����G���u?���=fǽ6�;���d��i��>��ѾEI?R���U兿T;2?|�5�`�>�2>�2;�+��3���4�=��g=�z ��|���J�K�C?|��������>��>�j�>�����s�=j,R���B>�Z>�1?�!{�{������^6���VY�̠��g>C��=	�>��v>�q����u�؆���V�>L?~�)�X�I>P�n>�f���SȾG���E>��>\q�?&�V���l?����4V������?KK�Q�E?Ŏ_������.���F�G�r��[�?s�<����cI�6�?�sn��De�MӃ���;�k��>K
� >�y��?>�q>Z����̾�9���vy���=3�����?iw�>ů+>n��>Zi?��#?oCK?y�ٿd势�Pa��.> gD?gD����M��GR?�)>
�t�5#�=Le���t}��׾�fR�&��=���>�Ob?�B�>�>��?g����Q�;|�Z�K�s?MՍ>c�V>��>]Zm=뤄>�B?��⽺g������,w��1����2��Ze?�g>[3�?� 6?C ���;>�t�?~J?��?>As?Os�>���=1�?I{7?k��>�
>���>�I,>HT?d��>�
? �?��>hϤ��K>;�0?~T�#Iܾdމ��,�A�b��{�T��?�pվ�%?�K�<*������0e��]ݾ1�/>O[������?�&p�*(����¾w^��T��p5?ϒx��F�{�>�j��Tc>k�q�U٣�y�? ��?vh�>Α��d䏿h-?�֩=ݖ�?��>�Y�?KKS?��?Ex=E��?i!�?�[>��t�s>��־��$��C���;?w��>�5�C^s?��i�2�>9bX=8��?4%���
?k`#?�Y�>�qʽ��
���`�4��v��"��>�㗿�V��'&|���?��㾷����&��?�8�ǵ>{��>7=�??�C?�g;���>��>����$�K��]�N>�$E���&�f����4>QH�>$��WJ��%�ʇ>���~'������/���k�i-a�L�������2��?g���^a�>��[?�?��6�O�U�̾N�d?�Z�'�O�"�>6]<<���mf�>���E|��UR��`������*��������f?��e�\�>������xs���z>��?����J�)��>���=�qᾠI����l=aj?.��>��5%�p���|ɘ���=Aid?C�Ǿ��?��>}-�����'?31-�;J>��3�;�8n��]&���Y��;�~�k?��?|�	���?.{���F���e�>8~�=H꒾Y�1>��=K�����>�����e���8�����.�?�V�Mʆ?��<���S>6eC�_?�걽W�:���~�`��>؊?��%?����'?a��Ŀ���?s���=T��>����ӫ�>G�ཬP?�=[&�`"���ɿ/[�*: ���濈+���?�Of��ľ�,1>#�?y2C>p����}�D�$�)�>d�C�V��>?�?��WM�I�\��/;�H�/��?G+�jξ�h�=�Y�>;���1j8?�lv�[�+<��C��.>F>�/���>9@��M?5E����?5�>�>��>Ɩ?VZ����<r=�?��%?�_�|�$�@qm>1���D�>����W�m�P��>+���<����f>�Zn>���������Z�>�q?a<�>M���q	�.׾��9��H�B��?��������d:���>(�cǨ>�;?��I?uq�O��MB��u�?cV� �k�Z>�?�>�Y+>'Z½|B?��>���� ?�&�>���W�����>����0?��پ�X�WЎ���?h����i=(��>F(?�d�>L�=��:?	%��1`���'�>D	�G�v?,>4s8�:�~=���?x��>M�->H#u?1�a��'�?,@���?�@>�^!?�Ɖ?>s�v���9 ?�8?��=r�=�ʰ�ֱR=VZc?���K! <��P<�@�?�ˊ�nN��Wr=�꾜�꾛ƴ�B�����>�<?�y���S�>�hP>�6=~�8?�=]?��?��
?����+�?���>xLR>����?/C�=}�ξ;dL?�[,>U�?H��>M�����������N?nCz>d�?��JG�>јn?ӊ�> �p�~4�x����-/?x0�?U��"��>Y��>�N�>��|=A�>�K��yt?,<��S�׾5�{�>F����*>�F��e�-�U*?L⏻Ѵ>�e��ʕ?\�� �M?����y^?�⽾r�8?Z�J�e�2>��>{���]kb�q�����=hR~=����p�־m򿛞�����8?=��h��>���?����TJ?2���'?��?@N?V6t��>q?�-6?%����V�?�h��V�>�n�!&i>�D��v���|��5
�8�ｨ>�$�۾?'l?�L��n�]�U��})$��?�:��pv��e�C3?VÅ�I�?�о��3#?d㲾� ��?��>�¿R��|�����+�>o�{?J�ʿ�(?���P�>}����z�=�o]?<��=�>��#K���P�J���?�_��w�>`��>�8�>j䝿�� �_�>��x=���>�𲿅d��(���^�^�?�����R��}ɯ>�?kI�n<�\���Lh>1q>����	�&��?뮎�fǽ��-��I���"4���F?Ӗ��>�>�_��ZD�GLw�'��>��>a|Ⱦs�a�"Ŀa>D�g�?��r.�78�u@�?��A���?�2Ͽߦ�>�ԟ�j,�?�����>�����U8?�?�>�s��߾�oz>[�>f�?�d;�&�?}���筆��� ?�p)=$K�>9=W�h�z<w§>�/���d>px�=�ԋ<�<?ƅj>�(���.���&�>�V?I�>��ȿ��=>� �> ��������w?�NL�ޗ�>����=�?C���q?�;,=�y�>�z� n~>V�C?�����n=-����?t��Q/=K/t�?�ֿ� ?X�?!L/��k�Ρ�?�T?�M>�Q���)�=��?�<?�3/�|�Y?���?P��?�f����<�QC>#�ʾj�����=d�ýjŜ���B��g=n�f�jd*?�>P�+����<o�>4���V?������q?�!o�Qi�>�JT�%�?>7�;�,����� 5?I
�I�>Q�S��D�>�[�=+��>V��k�|�
�?�F���BA�͛}?�	I���	?o�zu=ҫ�XZN?�c�<��H?9f?���=�e=���?H�>�>*\?�Ծ�JK?ӱZ�/l��,w==�H�>ss�>��۾ݬ?�	H?6�s�]�>C꥾���<:Gk>��?��¿���=8�?̈A?��ɽ��>��k����B�\����K?X�?���"%.�Y�k>V䉾�y?㏾Z|�8�>*��?�{k��vQ�H���4�?�X��`޾и�>���=�ͣ<��Qַ?�KF�=>$����{]?��������{�+E!?E�F����=�	�]��?�� �J��=�#?2��>򂿾���>*��>Oy�?7��>5W��>諭>�ߎ?]K�=�h!����?����5<�N��;��?��־�l�>��>��b?W�>�i�={ׂ���3?���6L�=��7>�m�Ȩ?������y�t�?.-��������Y��6�>�FE�Õ�q��a��I�������_��j^�����'L�lB���R?�L^����=��?�^��Ȁ?-�>
�<�?'���/�?[�쿠��?mr��u�?8aQ�8�?i-�>܍n?
"#�R�=,��>�׌?�u�����[�?J �?�˄�Ԣ۾�d�>w ?�s�=Ig�>~I>\[�>��>�%�c�= �7>��+?�H�=hw�u��N 2?�¾��L�>���%�>�1��	����q�%_;�Lހ?����}����;�ʐ��k
���6�,��>	A���Z��a<��/�>˞���zU�P>���.���Y�?g����)?-і���f�!>�?9�<��?��L>�eU�U�
����?�����$��ܴ�>mw��^��?\o��^�o�r��?ai�����:^ĿS"?�
>W}��}��� ��1KE����>�g����=��r��F+?�B��1���K?L?!(Ҿ���?�|=Hϱ>�U�?�^)?>O�=�(�>�I��G{?X�5�Dl��M����
?d��a���2?�	9?HT6��Zm>0�k=;�?e�>�F�>�����v>��0���ٿrx��0=�/��嘿���>"b'>rK{�B�-�J���.N���x]��`ʽ)�T�ɖ�>>ܾ9�H�<��k���t��m�>����eW��ؾE�d��r����9?9[M�Ϟ?f�]?5
N?A!�>�
�=�0$��<�>�uf>��?_�~���`�>�X?N�>�P+��p���>�k�K�p���?zj��G��=�_�>�G��<p�=A�����>�j�=�P��X��?�΅=�J�<Dr�J�Q?�̤<��������?��d>Y��̰>):P?c�?S��>��<?B�>!�>�̽>��>�M��T?��>D5�={���*����6>�t�>����>��`?�I��8�">)�:?S��>�f?b�����(�W��d%��a?[��=�½� ?;���?�,�OĖ����<	�D���>��߽1���ze=?��=�������#�M�J�CL?��y��bT�ǵf�k��?�(��cz�Tσ��G?�\|�r��=(�*���1? G?�X?��A�"�?�K<�O>�q�>D�	?�Ӽ6�?�u�>V 8�>�>g#��i���>��E��ώ=k�K>�)>[�>Ig\?_6?<>�;�ؽ�ܗ>��X?ne�>&+��$ҳ�}��V���6�=G���֮�n�F�`��>�Ĺ=�*G�"ú>
ِ>%g<���������?��?��5?-�>�^#?x�)�9Y�>d�j�>(�>�ﾭ�B��$�>�2�=���@/�!�:?��`?	��Й>����*���U��O�Ⱦ�j����=B�v>���Z��OǙ���Q�:�3�Ў��a��✾�9{�X?}P]��|�.hb���$?d>����="�nt=�f�� ��W����ry?�,�>��߾�K���<?�ѯ��#����>��
=5c>c�
<{���>MH?�]v?���>���ӵ�n��m�s.?e�ϼo1�< �=o�c��=Gx>[��}�U��e�	����1���=N����6���>�^?q�?�Ұ=g��>�TB��+���L�[f>�<E=��>#6�7'�o�>�15��E��<">��f>��-�h�r�c>$S%�iH�bl��X�>\J@�����C���B���e>6�?��=Hc0?5��>�@e�]v�?):#�|"�>��>�^R>�N�ԡվR��B��e�T\?k,�ެ������֚�K
�=�Z=YH7?�㶾���| h�C�?Ժ'�����!?�=�?��q�i�=��<�=�|�cA$�u.^�|��=^����n/���[<a�Y>}J��T� ϓ��M1?��}��ja����B�G��#?wܪ�4�����>:�p?��>�ي�Z��>��?�wH�b���]>nQ|�6��>=Es���>�� ��lX�$Q�>#���M��՜�R[�?~�>�Ύ������h>�
�=t�?K?�}�?�E�L�|<�z>�W���������>�lӼ�>)>�`=�#o?�I�=���t\�>�L�� `�>h���&���s{��u׾�:Ⱦ5X?��9>|�(�^���1�>�f�>� ??2�9�D�E�!�н�I���B��I�>����Jkf�$�>�G<�ؾϳe���>)�=`2.�B<���?Ǿ3�+>.�?n��>��5?��<k��=�&�0�.�`�?�J?�l>�uv���s�u�ؽ�GP?�?N��w�P>�Lx?S��>��9��>�L�>��<?����N>�g���X?L�U>�fG���`?L-_?3�����e���?}l*>
�n<�q<�;4>���fe?)�{>�]�>?�;?�G�>�X����<�^�?i;(�t��nQ'?}���N���n
>N@�>�0�?_ӱ�y�</g�>k`��<�>����KU>Ϙ�>hc =eo?7��aW��8��kD>kh�>h�>!�g>���>�Aܽ��4?�ͯ=��%�ȋt?��G��N����?:U?���>�?�oi�
����1�����:��(p>*;��+�<`E�c\)���=>��>q[p��2�N�!�-)Ѿ?=�� ��o3Ͼ�G�>��?� ?�Ҁ�*�@�,�?��?��<B ��
���+�����}�&��ߩ��(�=��)�
�Ü��]S�v0x���<|���'�<�7��Y�b�#���?9�J���?�x��#�=��>�"�u/�����(��>7�l���}s��3w�>����DN�9����>P���=P8�W�O���������=!L��{�#�r���dK��=[$�V��>y>�>�$>O�۾g�O�Z��H��='�!�q�>͢�<�e
���>HR��O������=�R��[B��0>�¾�ߦ�3]�?����N>]O"��;����]^a��"�=�K*="�K>4����>��>/� �@[<,wh?��>[�?)���	V>��-?Þ>耟��}t>O�?���=Ϛ��~Z?SA?�F`�r�>V���#��ҩ�r-~�13����>���=����AO�p8���>Pm��"�V>��Ǿ�E��`_?i��b��=�m	?�_A>f����%l�pP�=t&�>d	E��O�LE>f�ϾL�ܽվb���$>�@?~ֿ�u�T<���=���N
�ʄ>Z�j=c!���U������/>��*�>�.@��'�H)��E����d�0��=%�>??���t�G�"Ɋ?���>�y�=N�=�����;�?y>޽w�`�p� ����>��;����>��#?8s�>0�qp�?.&�>C3�:�?,v��K1?$N>�Ȣ�N~>Dw{���3���7�C�=@��>y�>ۗ��Q���<��9��?����o��n�>�G�>pXZ�k���D?9�>az�)�w����>�T"?�<h3��/'�� <�+"Y���b�R�>�i�>y�m>]��V�g<}(?�����A>��>�n�=>����?/�#<�c,�>���2O��� U>X���6�=������(>���>w �>:���9��q�?X�8>N���$����Ⱦ�'����?���3�$��>�5?�:m>��>@��>�)*?R�>º?`�>S���7�о���=��\?|�>|>?����Eq>n�?�#�=.��>�=���3>��c�I=�>\��u�Q?�S1?�q��SF��|*�=!2%?� >�Z�S�=���딤�p���"�$� ��ZJ?���������B��,�?�b���R�h7�>��I?����RX�4���Q�G?� -��X)�UR??��3�?�SI>ξb?��#?��c�C�b?��;?��>iC??���׾��=�I��7�>?�g>� >�]q>�;>�a��cg?p/߽�L���$?�a6��0�< ?Z�j?�`6?����/�=�>�H�� ��媽���>3虼UO.>V��>N�>��=ɐ�<j =�#?Cښ���>��־�l���R����Qk��f>U��<�����=CA?���¼���> w��H[>�DX�&���'��`����@�l��\;��g=~��p��K����(�nH?[�X��v��m=���gDɾ�:p>��=;mپ�g���/=P��>ן"��H2�מ�>�:>C��_�)?�!u>�4o?�`���>��b�*j��(�>g�̾&�>�� ��?��+=�Q?�D{?�H�>Z8J�Yρ����1(��&)>�񯾕$���ǁ��O�ı���P>��J�쒞<�~>��h�ߪ>vrb>QC�k_O��� ��>�䁽r��թ��8���N��We>@!6�pP��_�=��L��g����?�I���}m� �����=����bj�>��>?D[���|���]��ȯ?�x�]�y�mhl��Z�><��>��<���=��>]�?!���p�ʷ��[�9=��ʾ���fͯ���> a�qYS���Y�6Z��c?"��T�<���>+p�>	����|E?xڿ>ݟJ>@��<��{>n}?f8&?1:H>��@���>r���0̾��]�Z8�>���=в�<<�=�"��+^?y�9?� P�ɱV?��D?x�?�R|��oZ�K�ž��D�V�5�x��>���Aq-��-��<����9'�>~}��~9��ٽi�O�s��t�?f0��>(��>�����ELd���$�"	��v�>۟z?
���h��D��=v�
>���=������y�>5�=�I��哿�m�i�-)\>�㾾ӧ��-x�i�V?���>\4�=2�_��農u��� �3w�����I"�>�?�pO��?�.�>?Z_���A�kX%?װ����=�������S���5>���0��>�>���Ү{?Qe>���>T��>�A�>�=3?>I5?���}��>��3?3F�>��>����s�@?���>�d�<c��=FՏ?�?/?$=B�>}�6��뽵�<?]9?A�3����nF�G�ƾm@������\�?׉>��>�� ?���!�=}�?��	����g0�v�7�?�->ct�=|PO���J?��<6��?�A?�;�#A�<S��>3����O?�xr�F3��yH�eu=@派)���ھ��>�s�ޠ�?j��>{&?$��$"��P�>���?֌4��c���?�p�>_���X�>{�
���,?*�f� ���.?��F��1��Q?.��>Xy����<\\?F:?��"��C����S'��x�:�&:��JM=Z{�k+���c������J&��A��")�>M�Ӿ�߾8��ց�<�?MB�>8F?/p��B����=�m"�>�>��o���T�C �=9��>�DӾ�?�P�Ѿ ?�7?��m�~�=TL*?H�澁���������R	 >豄>�d���?��9?�)�B(�؉�fj����<F���?çp�{ĥ�}�?��Y>I�V���h<��F>G���'��u�Ǿ$�&��O\?�J�}龽��>⨥>��?ۆ#? |/?!-�=��>N�=���ZP��H�?��>�_>�}Ҿ����h���~$�1�����6?��~�x�>��?��A��!����>#�K_�!�`�3�z���u>0�G:)dﾷ�1?�$�?��?(n=�eh?��'�1褿MM?� ]?�����b�Z�}��J/�l�~�#�"�b8���>��<>���=uY�v��>%?��	� ��	e>���tP����qĒ�B��>��>��5>+e%?�Ⱦv��>n�;5D4�9Rh�ݴ�>~}��iɠ>�i>��b��k��5�> _�>�뾉">��������C\>3�
>$r=Rp��,��?S�?�t��+�9���A>��?G�\?j�<��	���>]aK��ټ=vG�r6���=�!��z?�c>����%Y���N��Pɼ�ȗ#���꽾���|E�	y�?J�D������\�>Z8�;1h=�dw?=���2W�>��G>�?޳��|�>&ҽ�sC?
, �:����_/?�g?�7��Bɔ�-�����A>�خ>��t;U�_�(>5MO?�����}?	<���<a>�6־<��vQP�	�F�l�=��=�Q;?%�?�Um�>�V?�̃?�׾��4>��ֽ�>n���e?�#b���?nʘ=��M���R?-=>�m6���=.��>((�>q���� �@�V�H�y>�QS��(y�薾����=[@�����>����O"��8P>��>�A:�H����j
����>��(?���>n�N?PJ����H;:Ri��)?ܖ\?"��q̾���=R��=i��>UW%?�@� H�>��<�.��4t�>�V/>���?s㾉�Ծx�C?l�>$���B��N0?�� ?i��>�Ӿ26�>�^�>ӟx>��J���`�#~�=����=�0?���њ� �>o�L>�3?���>���>�v[�3��d��`��>��>s˚?���>}��>��a? ヾ �C?%���Q9�+�� ?�+=�L��}ę��-�r,�*8m>��?5RB� ��ER?��>|4�>i5����>�y�>�W�=ơ*�S��>l�>m��&!d>��>� �u�/?�0?w�#�MI-��$�Ů>C7n���{��/�U#�>����}.�]��>`g��(j:�?K>�q�<z��?Ƶ>Y���N�(�� �>�?��4?̵���=d�O>��۾.�������b��dEоd�|��S
>���>E�����i�	��=JJ�>�?�Խ�̼�q�ʽ��>5E����?n��>�v������B3��>�2�>�q�a����9]�Ϸ5>��"�VN*����jt?,����]�}��4O׾%��e����/X��c��@�?��>�Y�?)���`J?|�1>���>�>ʾb�G>j��$mľ�k���=�]"?��͘пS>��>mH?h X� z����,�t�>�wj�6�G��I�jp�>�b�>���>[����>�P����>��=�<���������$u>�E>�+��*?zV����>�.�y=�Ț?:{���Q��=�K�>�j�����>Ӿ�>Q;���=�]O�-R9�9g�>R�i?ݝ3�����]z?%_-��LZ;B�=��9�L.�>0f�����u�T�o����%�`w*=
�<�v�=w<?Z��>�ߧ�+Ǿ�7L?���>J�ؾi��.��>q�3�e�߽C8׾��?
z�>�ߩ?٠N�-�>��,>�cT����>��>��=����NUm��?����>{��ߓG�5I?���?XR�=�4�>C�/?ڧ���[?�ѥ>�g>����&�> ��VC���=��R����=wFz�i�y�u�>��!?N�=s�?Z�W?��:��=)1C>o �=7�>��������;�:=Ҏվ��p�����?D�?��8�UY���xw?���>�c�=�k�<t�?�:?U�?��π�>)2?2�?��ؾK)�>���>!�i���h�RN`??՝���9?����Z[�Iȇ<9>lɹ��>��>k쀾f?;���Qd2=3�>W�&?T��ͯ/����>���>���Z�8_�>��>��>��V�v}?��E?tF>N��<�G1��5�?ت�Lc���??��˺ 
9�W�����>������E?�>[�/?��.�t�>����-#?��ּԫ��͸>�ށ?L�?6d�>��>��V>���>Mp	>и�?���=�Rf���5?�s�, 9?���>��"�
s��<�ǾPӠ>b��;�ĵ�(� �����z�-�1L��є�6�?�?ǈC�TоD��>z_�=��.?[d���>�闼O��>�|��#>�y'�|�>r��.��?^Z�>�5�>�"�D.�>���>a�=��<�?->�#N?ݵK�d|���;�>Sv_>K7��,��<N�3���>mS�AF�~q?�-�>X8>��=wT?�{�>m|�d�=�{X?��6?�x�q@ ��<��P�> p4���E�T#?o%r?F��G���I�>��?D!S�Q�֊>�eh>�����~>S�>�8i�K�S?�=�>h�9�l����F<�۽_A9���7��=����>E_�g)�^阽Q*�����=��5��/��"*y?]5��ܕ��p��==�-?8Z����>�3_��$>����"�>����oʾ���#�3}&=g~W?HFվ���Z�?�"?k����Ǝ>}�G=)e;?;�^��G��`?�	�=���=e����)?N'!?q�>N�p�	��*o?n��>�U��W�����Yy��Ԃ轶Y-�O�E?TO��\P��n5�Dg��ρ�(�4��WԾ,c>�ǖ��h ����x?�=��?��>�r�
G5?�:?���t�Mg=J��=�uо�?G���8���>6Eڽ���Ͼ \���C)?���=h��k:������΅�>��=kV>� 7�<�i?��U�~�	>�+4��	?��72z�h������T>���S޾�����j�>��m��k(�7�	?Җ�>O�|���\�ѻ�>�O��s!��kG�?"?,�����p>_0'?A;{=5"�>�x
�&�=ŕ�>[Ͼ����t��Z>>bD�[�b�Ԉ?�v?'������i\>Zy?#�>�v>D(�Wd	?f�����~�Ѿ@�%?K��\�l�?m��� g���b���N��M��>��4���ؾK��V?�w���%���0��s��a���裾���=\SE>�A���ez�8�:��!�>�>h�?��=�	?��2?~Y�=�6�;��?O�!>��=�[��
�<���>YQv?L��<��=�3þ�[>u������>�`��G�!?#�?+�Ҽ���='��D���QN���ȾL�����<��=l<���ֿ e<�.X> ;T>�G��9����>Ob�>��?�&�>Sг>��}=/'?I{�>|h?�:�>Ҭ�kV�7�x?�E?!�*?��r����>�i�>΋�>^��冾@��?Unt?�����h���C�x'��}R�������w">�+�?h��>�+?��6>7~:�,����Z�>�x�i�h�wz�g���(��=��Q>�_f>��;lR0��?3�i?5z��:h5�[þO#?{�r?�[\�xu��C+ ���>���=�����l�r�>�8	>���?�آ>7p?�4=�>#�,>U�>١l�{��a~t>R��>Q��>����=�Ⱦ��p���!����>�r?���U�ϾoH�>-2?���>�p���I=�G����Ն����	Nξx�ҾVɉ�����~e��M�,�>���_	�����!rt?^"?��-=��w�s�>Hx�?�Po?(��=���/���}c���,ؾ�ߚ;�[��i:7���ھ>p�>^�L�@����<>5��>P�	�MQz�-��;׾Or���]�&�}t�� )�[]�����>�&�L������������A�đ�<c]�>��پ�'�����Z�K>E����({���L��5?k��>p��Ζ���
�=�*$?�c�>_\D�����'?���>�Nd�ZZھ��}>p0?��d?��ݽ��?���ܾ	������P�4b�Hz�Y��>L�S?�C� �?/)�=1V���D��2M>�z�=�2\�㻸��3��>��>�*�>��>5�?�x�=��=��k?\׾������>���>]M�=ee��9{��$��>�>o�F=̨.�.7��~�>-`J�շ۾�y�>�"�>��u
���;�E�>o�=���`�> ?r�>�{��@�>i3�>"R�>�B�>������;n�=ukL>b����[���k�)�x������ؽq�a�B�n=kS�s4>�%?�w�?���t�>��>�o?��-�c���*��=��?��E�Ҿ<׃�L>z?����Y����r=�Ed�<c�6��a��`ͻn��[����Ͼ��$�%R��
%� �.�j��> �;?�?l���!>
*���b��λ>��Y>�Ҍ�8�T<�Z�?�>�P��a���L>!6�=���U��Y�=�_�>�v@>D���Ru1>b��[j5?����'|�B3>6·?.�Ͻ��W�+6�>[L�>'Z�d�z�+s��lAL��yv�<�ɼ]�X>�]n���=��z?�}��5�8�5\�PÙ>�>W+þ뱒���0�V��=�[��I�~~?�Q?	�!��7�iU��(>K叾���� ����OE��Tپgm+=R޽�8B��\=���>�})��/
���$�uA?�t>��>�I�>��>s��>`�!� ?�R�p�f��Z ��� ����>�g?R붾ƕ��B �Nq?��c?���3=Y�3<�>�?)?�?)�
�A ?ي??3Pb=���6�?�7
?F)X?��C�GA�oY>�R�?��z��N�$TϾJ�V>iоT�̾�Tf?��>��>9ʅ=����b�?(��>4�>W?@T���x�LoN>�9�?��n?�}�'�9?մ�?��C��#[>A��[�p>�s�?�E>i9پ}L��_�,�ԋ�U[���:2���w� G��5?l��>�}�=��=�Eo?ו�>�>�R�XR���>1�?B#����� �*�Qe�<�y5>4�	�_�B�VE�=X>�{��Q��h�۽�|>IN>>J�C=h5��#ei>vA?�E�>�,=FF�&�E>^Ă�l	M=��>#'>�v>�6���63>s?+�n=o��~c>93��������̾XNl��S��o!���[���8>�6>*����O���O!?�lz?a�>ڑ�=����M��v�?{f�>Cq>�����:���>��$0����ݽ36�;��:�	�F��>uӃ?��ﾍܖ��n��d ? ���ב<����yǾ�Z��/)���*�?[�=~�R?��>J�<�:���,>�rv?b �?��N��%�=t`�r��U�b��J�pX�=�*=
޾��=}�0?\���l���2�#<\��I>c��>������\R��c ?�cʾ���E�5?�q���Hݾ�� <�B�$�C?D ?���:OI�����L�>>�	�?��'�{�5>�Ž�E>�(]���>��>u�=�(����>��?���>���!$�=$�C=-3����pX�� ?^\��'�>� F���=�̗Ѿ�P^��Cƾ�c=��N��L׾�a�>ym�>�`*?��(?�n1>�E�����ح?Y�%���\���9>�*�=��>����
���>�)2?ؽo?8��k��E2<sk;��IǾwj>��������Q�=?��8�	�|�=4��>��3�>��>�6y>�6�>����7]���?�n�?t������C ݾ&�?a4�u�������s�s��?��>�� >�Sɽ��>��ľX�`?�����e��Gž�ɧ���ܾ����W��q�I�+��<���>>"?n;>tAC�`�>��t>��r?7�Ǿ�
ѾM9>���?mx��;���T	���?�Y뾐�=H�8>�>
�:��{�>�/��_{�>w2�ՀW��d������gy��!��"�t����O�>���s�>ص�>���=�i(�!����>�ћ�l#D�;(>-!�=��>\/�>����D�d>�tO>�R�4w2��lG�-��>���>e�������>�=t�>�\�>��t>���>�p?�\�>�c�>X�	>�>g� ? ;@?�윾Vv?y�Z��8�>�w?W�?��?�i?�=?����=}�A��9?>�>�Q �����>���>�Q >_v&��������q�=�{���B!���z�e�S���զ?Iu?G1>7�8�:��Z?&�?<�׾�\i�drC���?��+<^��4쬾��>�"�2ؚ?���>�?r�l�<�YW?�?p-���_輟F�+�3>� 	��\����!�*'�<��>�o�=I�����w>�PC?#�?�>�����Z�ch�>�z�?gzҾ��ž-������/��,c=��~>ҡw���?���>?/K`��'��;�5��>���>�޽3a����%n������zE>�ﳾ-i��B��=G�uފ�J��P�G�<B�=ĭ�=��3S�c�=�x>�T)>=h�*EG�U�3���j�T�p�������k��o=T�F�����< @�9`ݾ'{���:(?�>C�7@]�9�U�SQ(�L�>)v�>�$T=_a���b>UM�?E��>��@>�� �8�n���'��~��<�ǽ> j>?8���9��#�5���>��[?[餾&���1>�9?T��=�G*����=�?�7)�p�3��%���u>(ll�\a�R5�\�#�>�>�4����ۿ	�>��>�Mz>9$ż>�>� ������sF=�ڨ=I�_��㙾Pb���
�=�X<�C��� ��+r����>=��=x���d6�@G��H��;��=�>�� 7��Y����=q��>�fx���9�zj5?h5�:��>���=��A=�;2>B��`��9>��r=%��=0	���X��mX>��Z>��>��{��'>T<'?ZP�>*�=��?A�>=+�>h
�?ڵ�>y�4�U?(��=��>>���rI�t�P>� L?Fl??x�^�2�� S�>e[C��34?~?���>��#��Ү����=;��>t>�\@��*}�e�_?͏>��0>�˾�-�;Թ��%�	~�������6����������6?ߣ�>�)�`	��1>X/�>� f>�>T�V�n��B����=9y~�ʞ�>'����<�ʬ>y��>�0B?Q� ���Ŀ��?�'�?�`X?7��>F�T�u��>_�Ⱦo�F>�R�!Q?��(?EȾ=u�2��Є!�}�A?NK{�3V��a��t�����>���=�w��e>���=���#X(�W�<��>�?��fc�=�=
�z>����ξ�����+>�밻^ =7�2?"6�>8Ƚ E=���?�b>�3>Eg=�^s��ȳ=GҼ�x4>�3�>+���O��)�>,Be>=��=����7>b!��=>�5>���>��>�w��MN�Xx����ɐ7>4��=×��?�>=�=<F�c���ƽ���>���Ȓ=1�M>7�C>�>����_��$y���?�>��>M��>}���j��3%����>Iw���u&>:�>�3?v�O�����j��>��x>� �>O>�M?�9c=�,�˩=;-AR>5�>��!��#>�?>	�R;f�H��A�=�M�zB��&�>\��Z��=7>=��h>��潸}Q�>�v>D?�>8k>v�^ɫ�ʚþ�<����=����2�3�Z�Ca?�t�<m�'�	��7�?��>��n����d��><#�>W�>tk���>O0�}�i߭�3�V>�= ʽ��F���>(�5$���p�X��>�>��k=��>'��^¾���E�!Kn��d�;�`W>C饾Ӷ >�ýAǎ��G;���5ځ>7�<7��2g?i��}ξ�}!�"��>��J�#�����5�>ޘB�N����*�mK�>���>ms;�D���̽x��=C��>f�=����=?&!���������Lv>i_�>k��>Op>L�߾b��M��Y׾��7>��ڼxL�+?>>���=��� Y ;ݗl>����х<�)t>�X�>ݑ�>\�˽U+�<�a�<��=`n>�?�;ݽ�%��׭��#�=[D1>�����1��~��y>C�=�ѽ�B>��>Mm�= 쌾�ɰ>�u��*>9�ѽ��y>%p�<� ݾ�����~޽��>j��>/?�;�>���Qg�>	�>-G3�4�>��-=ݍ�=����V�>ZIt>���>������R��aiо�8O��0���>�V�>�ƫ<����t�7�sB�<�k?��=�%�[>�>���>��3�׾e�v=�D�y����L�fU=>�̼ȣ�=��0��Hʄ=Pև���;4���bvn>t��=��(n�9>�_��K���s���B;�$�>��>l7�>��&���m>�,'>dQ�=�G����=Nt��K�1��ϲ��\-=E�<�g��n��>߄A�'F����<d��>
�m�Bk��L�M��>5�=+��>���>Hy�>��\=q-�=F��[Ѿ79>4�x>7:?I�ž�2��ޝ���
>葞�ޭ�_C>�<S]w��} �C�;=
7�=�T���	����M>nW���N�x�>m�3>S�E��AѾ�� ��֙�9�F��ܰ=4dL���x��D�>b.��YT8=�N�UT�>��>l吾I˫�|ѥ=�I�>o%�>�$?�]�>Dͅ�����"Ѿo��V�=gY>���R��u[���(�>��>d�½��n�܄C=��E<"�	�7���	?�ͥ>Ϯ��1ؾ��j��c>c�>a�Ⱦ/�<���<��=� ��>��>�U�>|�ɼ�̾�Ҿ&�&�<j�>F�K>T&���?�>\����_�>&J�<���U�^>(b�=t6Q>��H>z���z��>x��>�`>�|>�Wf<R�A�^�`>�;=�m>%C>Q
�>� ���������f���D�,�x>�Y>��N��p}�+��ׯ>�z>N�q��� =P�=���I2���]���4H>['�=p,g>g���!B��9�>�M�>�8�=+ž��]�m6K><83���;=��=r�>�ܤ>sMg��0��1^b>n��=}��=kJ��_;�>ԙ=�>��5���>�Є>[2>�4$��W�<=jF����z�žJֽV���^����:�7�!��M�=��I>㙞�+P��~̽��=/�_�b��S��ě<^�b>�=��>'0���m��蒼��'��=�?ؽTƖ>�%�p�¾�A��wZ�����n��<��>�k ?��T�����&�9@Ѿ�ζ>����M�?��	:�=?zt>��>}%�h�J>X+�=�R ��#�D���ڂ�$Ƚ�9V�(�Y(�>ܹ�=Zǽ�����ν���1�1��������=���=?��<#2'��s>�ќ>[��>뿇�vj5�B�>�h�q߼��(�k#9�;��㢣��!��w��Ⱦ+>?R�޾ޝ�����<��>��z>�;>�8߾୐>�G�\����Hm�ب�>V�>ݱ�<�[�=�.�j��=�>�
�l�»��H����6�2���=��>�	�>���a`)�J=�� v����0�?��>��>���=��>�C�<�x=ib�F*?��cٖ�����k��=d�>�8�=1>_��>�/>I(H<����F��>��h>�gڼ��������Y\F>D[}��@Q<��R>}�b>t�=�o����(��:6��g�>I�9?�L>||���z齖*�>��<|�%�Rΐ�H�>5O<l���g��5��D���y��>8�1>�1G>`槾��>��d>� �5��e��=�A�>#V=.-��,�=c�(�e��*۟���־�-�>���>3o>>�侁�s���
>E�?ԝ��Z��=n�^>�Ђ>����K���܆>1��>���w�=�#�>.�0=}-)��[�O"ļ�i��r��=U3[>,�>1̹=��N�B�z����Ys�7��>��a>i,3=���>3�=�SR=|5̾�F?��;���E�Cĉ����=tH>����Ĥ=���>��i>N[>��+����=7M�:��
���:�-OӼ��W=^�s�N����4��7�>=�2>맕>`��>,ۮ>^I>��=�9�>gI)�O򩽴�1>QZB>8��>���:�Ć>AbA=�X=��=JKs>DW�����7>���>�
���4�Z���Ot>�B�5��WN���;��;`M��	���㾤�þcG�*�>`�o>T�>�겾Y0K�%tӽ\m�>{Wu�>,M>�L�>]��>�ܱ��6�{߄�q��=���#=��>j�=[�*���½`�L>��P� �:>a�>>���>�+]>����x}��F�������k;�'�Y>[�>�}���ڒ�v-�@D�>CL>J�E�n��=�Ԛ;H3<y�v��O���M>w8!>�����C(�>���3�����܈>#��0�t�䙛>xmK�2��� ��cK����.�8���f>��a�������>�T�>��=NV���b�Ni>���p���+��>-ke=���n��V��eCR�l�½*P;��_i���=�4��A8m<弣��c>Vur<���]h@������9>��K=dSϽW�߽�T^;�u$�����t
���i>�Ӂ�E�6��7�=����<~��� ��H���^>���	L ���c>P��>V��=E�����w� �>��7>�+��<=��>t�>��ľRQ�}��=`�=8�@>�a��b�`�q�t>寗>� >d<������gc>���b�>��S=e�v>�r>��i�BR�DӢ=G�9�r*`�7N�>��&>A�������������>:cѽѦI���[=�l>�	W=�x;�N�eȮ�"�>Yh��_՘>��t�!�#�ݾ��ͪC?8�+�«�=f���1>��A��o�g��=��>�k�>����X���r>U�>=1>)�F��"!��0>��ѽx$"��WS�s��>{��> �=�e�<���>� �O�;�
�>�k�:f,1>�>x�|>�Φ>����og���s��.>�+�>�0�=�>?���חl��6����>;�r>�b[>Q+��j��>H�:�G;�D��V�>��>%�ͽ�dľ�m�>'Wܾ�=�A���>&��=۴ͽ-��lr�>#9�L�齲6����>���>U���ֺ�B��"N�c�J�Өi��?f���	c;��q�ʭ>��~>��> vJ����>_\>��;>Q���x�>S�?�j�=8�
>��Ծe�˼WW/�vr�>R^��s���nŽ>�@־�c��x��c��>
> vt?�5>j�=9��?�49>��< ����!?�D��9^�^\#��l�?wS�yL}�(���ٺ~p<�r>��H�P�&�_�>!?��N>�ŗ>�Ό>��r<Nџ>���>DM#?��=�$ ?"⎾�>>�Ư>V�=�a?�0I?ςT?���>7(Ӿ~�������R>G�&��A!��֠���+��K+��)<?U�>���<�I?��=�$�/�M>�� <�Qm>�.�\�>�?��������7>>��>��t��z>Ǻq>z��s;�=�T�>-_O?�Ҹ�-iN>ſ�=`^�>@�}=��[��D辬� >n'�=|~?��?��>R��?=�>���>+���-	���>�];3��>�N>9 þ{����>_'�={�0>�C>��g���=0>9?3'H?�|�>ZƉ���T>}>�������̽��N�\���!�5����<12��6K��HϽ:�Ӿ��Q�� Ǿ4��}��=��������Z?��>�t?�_>�k���m��MG�=������?��>e�l���l���?��½�҂>��򾧊>?2�>��{=���&�?h�'��$�
����i^нV%���ʹ>�<��t�Q��C�����<�)�Mڊ�n�q=7g	���=�=�>w�޽�(����>nľ����N��j�>����sG���(�� 7?U��Ta���>t�o?u�����0~��`"K���<?ff�>�Ј>\8���d�;o�����a�M��O���w��6����ᶳ>4e�>1e>���>_NG��+�=��4������M�2%����`�;?��ž8�����>��~=eN5?��H?-e^>0�Q?��ݽ�j�U����>y��>>����=H���&O��*��s�����Et����Ӭ�>\�R��+A�t�Ɯҽ��Q������g�=�W>�3?��1>��D>��?���H⏽;yb�(�%?�"�>U(?z(x�`�˾Y��>X�>�#��h#�4�H?ʬ��U&��Ҁo�WwQ<?	��g�Ͼ���>�B���2^�S��?Z��>�8�g�K�l{&>�뎽t����>/��J��> ��=�>���B�ƇF�l	��D����W�{N ?����
^�}!�>�N�>\:���A�>�)��k�=~<c?�;�>%>s�Ⱦ��&�Q}l><W�=Jo����5?���>����(�,�B���<�yŽ�h��r�7�M����P-���(?Mn�p���V�
�ƌ�>�zX>��/>@#>��?�k?0m�>�	>I��?���=� �>d\�=_�T=�ܬ>��x�>��z>zP?���>���X�����m�
`t=��<{�;��>?�t=j��.�$����!�*?���=A��týK"�=J"�Ј��荿y[�.���R.�j������aսݒ��;B��3��۾���\>�1>=>����Jf?s%�>��T>��?BJ�;�[��u>`%w�QϾ��pu,����>L�Q��yJ�y��>�g>bw�Cs.?C%�>��#?��>W։�%�4>{��=�.���|:>���>�V�=� n��5?pi-?��>��˾}�0?y�G���C>	@����̽�iv�p3e�[�]��K�>F�=���>Ut{����>+����FN?�?+�*?�t�?4��3��=�*d>lˌ?��\?��L>yy���P'����=e������>�t��1b=�%�;au���=�ʽ>�j���?�3��c��>�2�U�?��f?7T?GQ羊�6?sXt�_�>i���L>��;ӓ����">�bh��.����J4k>���2����D~"?����o�U>`$5>+چ��?3�-�:z���=��?oL�>�m�>��H��Y=x�k>�(1����=�=־�P��jK�Z)��xR�����$7��"8�"�*�2>=�K�ҽ��K>L�>�_�>�h߽��<��(?b�>N�O<HV�=�)���K�>��=w!�=��}��n��q��>x�.���ƾ���K�?��=�%�ƼS�����;?�@)�G��
ֈ�4.7=B�#�'�;�L>�;�<��>E�=�� ?����M?��!?�yW? �R'�b���*��Ğ�� (�~枾pL���N�<Mݯ>���>�5���b��?D�\=�$
����>J���GY�>�d^�x"�?*�?���r���Խ?���d>Ng5��r¾�ld��A9>�Xþ� �W?1��>t��V�y?#�?�)4�vw쾈��>�t>�b?��΋:?�E$<~Cu>'�Ҿ��������W��i>܍d�B�>���n*���#����+�u��ϾX�ܽ���>�+�����&��>�ܽYp5?�B�=b��>�]�<?�S�"I����^>�� �g��n~>% ��|�|R_����=d@��bm!?� �=��L=ŷ�>(C-��<������JD뻖�P���)�D?�C�᷼�f�;|N�>�>�ڽja�>��G���?Ҥn>�Pp>�%	�� 
�;2�F��>���g�?��������?l��>��x���&>^��>�>����1]<bgB��g�>�0�>����x�G��R�ƾ�x��z��Gj>Spk���L�W8c�A*�>=ђ>3�y����>/�U?D�>?�$��=�X���`�>��Ӿ/ӄ�����M�I?�Q��4� ?�1.���>QǾD�E�B�%>�>gf�:#I=�7��)��>��������?��>3_e�8��=������T�L����Q��<�=��>��>M*[=p`���'>v�����켵Ua�Jn?�?K���<�~=�m�t�&30=�=�l�z#?e��=��>>/�>�3A?E�?e�T?�\�Mt?Y�/>���.x ��"?f�m?9�þTI�>`�ľy{� ����3�k�=��9>����j�>��Ξ=��C?<ʚ�7]U=��F����>OU������������ؽ=���7�.~6=��k����=(F=!N�����O?���>Ty��[)�=�J�>@�;>��q�$�������'�>b�r<
k?Nu>�:s?s_Ѽ}U<?uZ�?��j>�e�(�>dE����;���>'�J��|�>unվ!��'����=�>t������>�r���{�>� �V?��]?��?�y�3`�>�F@��j�>^0}= F==����D����O�~>Mު���o>9��=��>��>��=�U<��{�>���>j�,��TS�~"?�>����Ҫ�>Is����C>F~��X�>��ѾhzX�#k�P ?ג?��{=H�þz����(��q�o�r��T�¿.���.>�L�>+0��V羛�>󔵽���?���>�8�=�����a�cA��O�������"o/����n�?+a?��+?�j������c�>_(�>}�A��)=��
?��>�;?������=��F?U�c?������.Ҷ<�'>XT�.�#�$�ϾJql>�>i�>6�½�m�����>����T>�+ʾrew?����RMs��6y�q�>�R���ZN>��ɾE��A�-?^|���"2?�c���M�:ꊾ	HT>_&Ҿ*�z�
2�����>94���4g=�e¾(K�Zi�aV?�k�?˃�=*�����=NQ�ޭ��0��=~4����>d�>f/����?_>y��̼�=�<+�Ͼ�Z�=�
��N�4u��>^&���4�M��:+�>%�l�&��>��Z>Z�>��7?m�D?��߽1��?��=�����5����>�3�)�K�;�>�E�^�����1��x��=;�?��>4���S?z�= >���sw`��f��c�Ǿ���d���U��O��n(���@��j�>.-�-3�0�E?fM��z�.X���{�=�����dC�U������?lR6��@>���
M�������>VA�$♾�g@>xT>�4?b���TYӽ����dŋ=]� ?"��>�{h�'���Ek��&��=Q�:���(?Ej��yN>�"i=�f���9>���C�>P���a �f�8����=Ch�>f��>���<V��.~�>�'m�h�	��
�T%>�G��=.Ϩ�U�c��P�=������K�G�ټ�3�>"x��+�>�3@�Ħ��˳>1x?�ؼ��@>#!?�F�>��V`�>�6?� ?Ds����>q�>K�>X������;���>�4�>%�k>҅8?=�4>��ݾaʾ�� G��g��@����>̎j=G��>*?bȘ>�*���Ͼ�k����w�Gҽ�]��÷��,�=��Z��� �<TH���꾹���>_ 7�ʰa��C��Ber>fb���Z<u+��͏=����������ޡ+>-Tu>�>|��>��y?xVX='j�������{>C6ӾD63�ٿ1��b�>q�ҽ:��=f�a��>-�����>�WU>^����=&����>��?�㤽��v>�$3?��z>���?u��֎��q�
��!ؾ\�ᾗ������N����>�q>�f	=�^�a��>5�=���,=m�����>�}U?��x�55�0�=o]3���>}O���i�>�e?}��IiP���>=�Ѿ-N߾WA3�t�"?���<�7�-A�@~>2�>b݅���sǾ�����T�<}�M�1��?������1i>7��~�t=�����ʾ��<����BϾJq�Z(�$ö���F�<i>�'�=�����`�Fc�>=b&�}Ԥ�|)o������= $������l<��K�����>�TI>@ɧ�h?Bq�=�?�����k�оηνVD�=	?�̽\<����>6W�>�z�: ӽ���C��=ɽ��r�=�h�>+*0>xPo�d�R>G5?Q��>�Ƥ>N�1?ww0=?/���/������+��Ͼ#���UO>���<œ���
�=���>OD��P�˽|�%>8h�>�����Ծ��<��(T>�1� ������>& ?z��>�ܟ=+ɽ=,Ud�O��>�m��2��+P��%W>X5 ?�T��.D?@7���J=9l��;%�8.��e���yS���+>?��7!<���>©9������=���?�Y%�^[�� >4�(?L�c�S��P�>U�>�jE>$�پp��8{��Q�M������l>=�>�b���2��:1>���!������|�b>Tp�>��
?����g���?��?[��+��<�ua?0��>.=��C�=��]�� >%�̽�J,��YǽL����?oR>��Ǿ5jr�Q_	?������z������a��?��s�TM>�գ�&�>��?�轾 �6��>��?g�);r���3?��>�;�K���^޼��X�;� �L;J��댽�*��K�=�j��{O�>��=��	>��=�QP�>7�P�Tv=:��� �:��g >���<��>�jپҁ��H9=��>4ܾW\�ˎ�=M{>A���}�!��>�2�>J�?xv>��`>��!���پ�G���� �X3Y=	��>A"}?��=9�>��!?��>�V���9�>��?� �=<�=�}����=	��>o���)�>p�>"X?�3��J��O&%>ձP?3w��n9�=�k�>%>�>��ɾ��{>�� Þ���4�6<��p��<~�I?F��>�I�>Ro�>�>i����^>��,?C�>��'?ٞ�>��Ľ-��>
n0�}m>�!>�k:>�^>�d�xҾ�P�͖��k���d�����1��J��>���>�ǾW�?>j�>0n�>!8������<W>�?w�����>���>��=n?�}1�/�����	�7��>O�
�ڦ0����y��>�>����ѽ��+���>P2��QKѽp�->k1n��ă>9B;__O��x��?4m>��=�^��>9#�>���>&Y;�F����p�TH�����Y'��I�4��5��	�~���(�V��>���>D׼�@>˕�>�D�>���B��;�����>	� ��!f>���>$I�>;�?����G�}����Ut�>5�`��0��1"�|'?
j�[�E�Vf��>S=?�w5�j낾�y��
5g���U>���>e<?d��*o?O���^5>��z�<��>l��>݉u����ϩ������R,���/h�[�>�ʮ>�K4�H�>è=��=:����]>X�ӽ��?b����8�>owX����>�b?�a�;I�X?;״�*���V��	���sP���"��O�>o,	��0M=���;�>��c֠>Ż>�6�X!�=D��>i��>�R����K>��9��d�=�P4��`~?x��>T���*����E��Y��e꾿�m��>!��
�>���>w�=p��>�S�>f�	>F�3�پk]����0�+oY��?��=��#>!6�>Xf�=��8�h-5���E>�x��%�`.��T�?qɱ>QG�=���=S-�>M�	?�~+>�\D=��l>V�>є��]�Z�N�1���=���;����/����\�=�-��� ��T�;�L<y�"?�
?�`�>��S����=4n=�����oܾ6�>(�����'���e�Z� �����w>&?q��>�4y�'&��;�o>{>�ξ��5?ҏ2=���
�6گ�5��h�����f�_��� ؾ��">ۻ8?U �;W���0>k�{?�Z���*��n�>���?�/���>��?k:�> 6�;h��v��H*��h����Ot>�<;?��O=l9�>��>^(C=o�����*�������{�2�6a�>�!��p�X�~3�>��L>s����i��t��>��>wK�)����i?��>��>�eǼ"bQ>��>.﷾*����>6�==/�=g���d9¾!��(y���A���>��)>�A?d&�=&7�>�o�>\���}>��I?�O�>�E>���j	�>e�;���>83�<�2�>�K?�ŝ=F,�>lϵ=�l>!��<��~>�� �I!���/�>u��>`�y��\>W��;��.��e�/=�D��G��q����:�;H�˾ЭC?��,�>�_�͒���"?Z,��f��a�E���?�}�7�
�>��L?TX�䰯>p�>�/輄=2�sa�>`&�>�_�X�=�&�>���>7��vMF=�D�� ��"�־���0ξP}�>C>�>.X��G?ު\>��>� ���@A��Q�>���>�����)�>���>�=�`׾�k�>�n ?��^�LsM�8�?��=c�+>��C���>ns�=�޾	�����5=(Y㽌]�>ͯ�>�J����^�w>��f���4� +T>&1�=|=��i�5�
oc>������n�l�u�n��K�=Y^��6{��<���B=�h>+w~=>� ?Fb��(�2>. ���*=��L��?Q��;�[�|�>jQ�>���g�A�5O;?�L�>��X����Y5 >F%�>�K��?���#	G�"((>�d��q��&5>�m����>�������Ư���/L?m|��p��>��S?o%	?[��`�{=Û?�R�>�؅>�)�>nu��/���l�>7�"��T���s��=��>���=ft~�ݐ���w>�+���@龓p�(ؤ>C�>��<L���Ȁ>>���]w��-��W� �'3>�����'u�1G�=������^�}h��خ��?ʾ���F�>��?�k����4�7"5? ��y�!�Pˣ�j�m=�Vݾ^5�>�4C�#l=���>�S�<�%��㌾a�?�N��	���BP�>j�f���Y!���>�G�=7>N�?\[?���>���>%J�>�W������!��`|ܾU��=�<������>튟>���<�-K>cj
?��??m��>�Ӄ��z��?�g+���6��pv>f�x>�e������{T?7�����׬־(e��~��>�XļMH�殻�봻��O�g|i��݀>/�#>����D˿�C?{����'��5j�a=�����i����y����ۡ�=Z{>AD�>��#?W��=�}#>���0v>�[�>4�?�=%j�>�(ѽ��o;���?lݼ>�"�?�5��=?��v��9�=���f�>�,��F�<太=��[?L��=�K�:�־��ľ��b>�↼�#5�ɰ/=�D)?V�l>F/>{ξJ>w�b�淌�䣿a�>r?��
�	G�=:��>�,>��y?�T��U�!>s�=d&�?�ߘ>���=hT�>�O�>i�=B�ý#R_>�D��E�0>�O>%��>��>Pt�>���>-I�>�g�=�8�]L��᫻��ྮUH>��>�@T�b�<8k}=����3��߀>S(�>�v�������=0�J��^��¾� �|����AK?�kD>�z�>9麻5�5?�=��>�޾�#?��0;�ȏ���	7���>2	�>�0>$<�?����׷��"ž��(?A��>�=�=���=�L2?Bs�=�b����� ��,R �����@�>���c'X�ΒX>a�?��>�pe>��->�P�=Y=N���3��䘾H���)��^@�>������ȁ"��o?�!>c�������s@Y>U��.�������?��ν���>$޾)��>�>i�J�Z��F>A0�>��I�����`��
�?��Q��nF��&S?�M����>�;3�>��ͽ�龡[�G�"1~����>�-�>���L>���>�!����<��<�������?�ҙ�r�˾�H��\>�\>^Pо�,н�%�>T�E>� u�qɾ���>`M���
�>ժ�����ֽq�˾��$>�w�<�'�=���>�'�?�i�=���>� >��>��U��7�w}��2���;��=Ao���ڄ��� =29v=~���}�>䕋>�<�A����ŕ=*1�>�����ž�<�\>;�?Qw�=Y�*?FWf�^q �޳���<��N>?+\<��=��� ?~<��T��p����>&>�in>�	!>G�>6��<r�&�pQ�v���:��5mA�c�4�$� �}E?�h�=W��=�>F����C���HZ?5�˾{}��{���>�3���?��Oþ��@>������(��U ���='�W��=1Kv�K��;+1�V$>Q��>W2�>���� �=�=?M+?
���C=��
�	�'?�Ⱦs���2E>�py<���>���>���>t�ԽAQ>7��b�>?h<���2���;>���>��>���>t���W�\0�>���VP9??;F�ɻR>"��>���>-��A8�=7n�>x��<�̞�o���ɼ�
>��W>{Ӿ�r�=e�%��3�>w9�T����0�ӯ$?�#��1��=d#�>���>��>M�L��Q=
C7���[�h���B#?����"���밽SW;?�ӵ���r�l>7�>k�<_�/=e��z�b��'�EN;G�='�$?��>�����jI>��?�=V���x���#C>����]�>�>,/�<*�&?-�����<���/�t���:�t��Lv޾q��=J�?�D>�Bn>R0�>
��9M���N�
�֛=ú�>�tk>Ht�;���?-��6L����> >X{~>26?�c�>ycB���>��>@?������*#�>�>���B/k<�Ҵ����>��4��[ >����B?�����G�=.�@���	���>�@�>��>j�?�"]�>�?>���f~?���=Q�I>��_>��:?���Y=>(���ȱ\>_��
Jc>G�u>E�t<�/?f�\>(�����>B��X<��� �T��������>�;?zڟ>�������b�>Adb����|����Uf=�ź>�g���ģ>��A>Nï>bc]>؉��O���1��>>*>�~���4^>c`>�*<�ʐ��*�U�Vb�>$���S�á`�@�����
S=	<�ue�>��>��:?�,Ҿ��?�j�>3��>+Q�6ɾ��]���f�܊=�./�X1v���=�mm��lm;�Qc>�,?�Gо�Y��y�=nD~=@���"�I62?��?��>"��>�-�>Ց�>�G ?30�)ƾ[���>�?3OԾ%-�=/BS����>z�= ���Q![��u�>�<���o��<_����l?��>sn�>x�\坾��ܽ�.���,žn��/�>�g?����B����4�U�Ž�y����<�xk>x�?by;d�����=X
��=��lG��>�?ɟ�>��ֽ�[�<��ݽ��?Ϡ�>�����;��N4��?F�\hо�t�>��>X>$������=�1��7f3?��!�>��a�-� >��h���0V���	?A�+����=B�(�ӽ>�S���w>2����sR��>�.1�F��(�?�K@?�;�2+?)�<�B�%�>�����Ѿ����u3
���>�D>?��v�/1`?dA��KeQ�ڸ��q�>�ҭ>�\*=#R�En�>.��>�	���.��Ïu>b$>�(*>g���Ҡ%�3f��:��J!���>D��>C��6�̾NG=��=�=���%(S�o$C>8ö�Np�>�=9<3(��՜�iq�>��?a]�>���=Ҝr=���]�ʾ���e�d�X[��%>�F'��>���t�=���k�>���<GZ?�PF>l��=&������RH$���,��? �sdF�M��>���>@��>�h¾8���V>�VH>���_�G>4��=�'?�p��A�>Mގ=�|z?!Ҿ�O?��	?y��=�6=I��=��>D�S����>.����I��{>������܄�^�5=j�v�:�>tӘ��&?��g�t��<�\���!�dA>��ؽX�!��F?���>�L�M�o9>��=���>�`1���?�!.�r
�=�����I͡�O���UF>�x>kx? u�>e��>*�>
m�>�7??9.�XdN?iJ�>q��\W��Jv!=��žJE�=�&?��ʾO�N?��>��>�m�W����]E�Po�1�>8%��>>��>�[<�P�?��t<�$>h������'y����k܇�VZ8�v1�������>3�f���>��9��FJ?�9��_=��u���?����������$>ذ:�����l>:�ھ���>a�>GqC>y�>�t[>�<�β>;��q��w��)�P�����#���g>F�?	�>�w���ؽ��=BuO��5 �+Dؼ��0>ek>�����(�>�y�>�u�>vG���
<�;�_v��o��4��?Td$>�?���=�>1���Cݾ���>A�x=I�Խ0x�>��6
�17��EG>���2���!}>S��>b=�=���%����V�>_�=� ݾ����btƾ�N��4d�,�z=h	�f��>��G��侕�Z�h&��΃�@���>�Xj>�(�>~���9�>h��>qA���� ��Iн���>HƁ���%������?-L�<�w�<5Te?�!�>@�˼c���-�>b�>�(e��<��==�v�>�%?� �=�>�y�>��?�0��U�=��׽��>6ȣ>�8��V|N�A�ʾg��>Õ�=p����_>��>���5A��Df��׍�>!��򲾃t����>1N������R�~#Y>Y'=O�R���(>1�?/��=~��=����)�B>2CX� �t�ݪ]�Zc-�m*s>��>gҹ>�:�6��=0�&�î><�Z���5�;��s^?v����>��
>��4>S��>�V �J���l���Wi�>(D{��~����=ƾ>b�C�AK?�݈��@?����]��d�?��o?�|?�9b<��#?z��;i����=��>��>��>Ү�>�O��#�7?�𜽯-�������?�F��ǜ����ާQ>�-����C	���
?n)>"�#>�{b�X�i>_���Ԟ��^���v�>
/�w���wξSզ>���V��FȽe
?,v�=ϕQ�4c(�U�>H�!�[(��a����M��P
��؟��PV�;�)?���>���>Wr���kѼ��=C��p�;>�->�.?S�V�������|>���V�=�{a�bh>����>�����K�>��q<4��>a'����r>l��R�=M#@>�C>�T]� "$>�@>_ɾ�t�o�J�	��=��O>�3�e ����>ə>�H��
Bf�Q�ž��>g�<d9>�4n>����I�"h�>狒>B!��￀�ec�>9�>�������=�w�>��>mk��Y8���	^�#�ɽB9>{�ټk��j�Y?���=Z���	g������-Z�������Q>`K�>េ�hʺ>��>�ྕ;��� �=<�>�#3>L�k� 2�=pC?�5�����Vu<�&�$��>X�>m��>�oq��L��/�&��}�>��0=\��:�νgI�>����h�g�.���>U<�=�?L���8pU? ([<�j��w�=J��>�:�=�i�=���⼦>�?�D'��B��	��=�=C>e"��7\�=V��{�׾h=�=�>�=�7J>]��>~�>S2���<��� �	�e����(�;����N@�E>ϼ�=!?Ba�$��o����=ts~�����h�2f�>��%�>.��<�?4Sо��^�FP|=�g�>|�5�d�l��r��;=�Ծ&��;�և�V?�)�;65�>U�==���>��a������4���Oʽ�Mo��=�>��g��7���?��=�87���r���e�`��>*pϾ��?�f��\Mɾ_��=���=iN��$�]��տ�=��=q�@���ѽ���>*����=U~�Mhþ�U>�=�=(;�>�\�����+� �=]A>���=o�=�K��28��F�t�K�5�S�@iB>��=�!�=c�>�$>���*:��'=�Nf>@+�h�����=[>�>����\0<=&�=j@>S�P>j.�r�?Q)�=�+���=ZU�>�;;���<J����*�=�1?z۾W�M>8����C>�K���A��0
p>�˙>G��<��u�=&�p�k�
���Ľ
��=%-?Z|�=(�.> ��>vF�>����Y�X>ʗj=�ҽ��a�X}�<�h�?ֈ>fʦ� �:>��>��U`�ѯ���:���b0��C�ٻ?��S> Ț��6����=Qq~=�-_>���N�>p�=���>)�;�!>:4��JO�>��E=�־�K#J>���>?ӾU��=���z>)*>�t��83�了;9����E�>$�8<�Y���X>Ј��q�5�<Q����t>�8�7�h>/���4{>�!>�:�>Vߖ�*O����u<��<����4z�`��=N�ԽK�>l���I���M����>��������s����]>Z��>iX�=O�=���>���;�녾KQ��þ[=�C�<���>�B���1�����>`
1>�9��tS�4���@=�p�`|��M�=��=%���pG��h�=ͱ�<��������!c<~�?>Pv������>���-4�A�=Lo<=Y[/�ra�>3%�>��F�K�삋>̆��xc�k(~��(G>c��>#��>�q|>�R�>^t���ͼ�%f��^����=M��>*�q���D�3�Ò=1�g>dL�=f�4�+)J>�PP;�A>�5'��*�>9�>�G ��u�����>Y�='X(>
�ϡ ���>�3����!?���Xo>�+8�ֿ9�2�>���Q��E��>D������=�I�>,���;�=����ܟ��C�>��i��+�>}�>�Qr=�N�>%{8?3��dSi�MG�6�>��>��;��1����`=d%�k-��򈾌��nᎾ��b>���>n�h�!���*S>B�=6��=_�>��ℽI}�>�>�^���t? f���=�v>�����b���>m>1Z�\A �5�	���0>����Ic��>t� �?>�־$o�=C��=�8R>�Eս���=�R>�"�>�}�=��>�k��8x>�"�>ґ�>g�ξ�����`�o�e<�Ժ��+�"�/�K@�=��m�ϵX>�p>k!����¾��P�Q��>�.z��엾:g
?H�m=_�Ľ�0T<�5���Ã�>u����;�'�=�M�1[=>S��M#��l�?0>�Y�=��>�"�=��e>�}Q�����`�d=.������=v�>�Hy����Z��=P�!;즣>����a�� �4>�-�=GJ#���=��徨f=�2B��	L�W'�>��2=R�����W��*���>Q���������?��=L���^!<e�>P���=(.j>�����>=+C�����8�=Vzg����-V�>���$t+;��_��%?T�
�5&��?uV��A~>wS�r+;��X:|=Z>�<T�f�=m���(?2q۽��>��¾M-%<�\�Z>��=��H�1v����=�c�%%�>"���sh>"}��Mh�+�_��ھ�:��H�>XȨ>�|�� ׶>K�:��-= �=+?^��=*����M���x>@� ?-��!��ĝ>Jy>�=E�Q�̍�>\>�Rl���[��8�=���>ۖ=����e�=R��>ʔ�+䔼��=�a�=��=)%}>7Ь��O�HCe>L�>w�u�mh>{���Cm=�)��言����Ք�G��>Nc��K�<K��)3�=���=4ش=�v���g�>�1q>�[>\n�qzN���Ⱦ5�@����8+�J� ?oP?����1���.>��V=M:>xH��|(�b��=��B>�m����>F��b��>YD>鋶���>s��=����82��-=Ps����>b����<=rq�I�W��Ks��䢾����"a�;$%>���<r��>g��=X�L>A�z����=!��>�-��'P����>˩�>�kW����Uɱ>��<��ѽ~=�$>��B>b�=W����<ut[=o�5��l��>�*8?���>;��=[(�>�yƾ�r?���m�>l��>>wU�S?->ꥅ�%M��顆>4[���ἛJ?uQ̾,z[=y]>A^�>R=/��^D��>�V����x�n>�h��iMb>Ay>�H�>`싾Z����ɾ��$>L9¾@�k�#��>�d�>��>K��_'g=��L���(?�m^=<>j0<�+��>ǝ���9���/ �})> �7=]�>p�E=�����D>N�'��=޻G��Ç�4	?�h!>�n��K�u����mŽ@F��􂚾JY>�u�>�d���2��� >��D>S��=���E�����>��>��F�v�?��ż�h�=�(��6p�ld>`��'�u�*j.���_��j����<s�x<AP->=����W(����>�<<UJ9��ͧ>��\��(���i�>��=�q����p���"[=��(=-V{�K0��>�C��X �[�U��)���Ѿ�=5>x9�[i��<Ս>eU��g���M䎾���>�j����^�c"E?gCŽ��޵���SJ��=�>�Ĵ�
���1�b�D�h=�f3�_������<ӣ�>�[8�W!����?�w�$�b�pO��C#?��o>D/X�i+����=/�*>_~>G�Z��[�>���=�-�>䫌�[�\>�	����M=��>�e����ɾœ>�X�=z�]�G������^]>�>�=Z��l?ý��>F�'�Dؖ<��ؽ�ߩ>ɸ�=^斾e:�>�H>i*�����n�U=�[.=Tb>H���/ʼ�_?�?q�۹�����'��o�>��O>���=�<
x�<!�Ǿo ?�g���I���v,���>Ǒ�>��6>�靾�1�>�Q�>{l��]ֽ,�>>��>`3�eI'���"��5�=�1�����*�ƽ�e�>ڎ�۴�=�o�=��>��?�8��0�>	}�>�Ҿb�>� 7>.і�`ـ>I�ؽmrN<4#0?�4��N>Ř�;��?�+�S��{)\�^[>0fq���=�߽.C�>��>��=��Լ]����W��	������}%?W����2����ֻHz�=񈄾V�H��d�R��=�[�=[.���/4�ڣ�=R0����=��Ҿ=�<��(�N�:��y�D^>�n>�����夾}-|>��	�=��=���:b����$>im">�D�=og�S��>ND@>=E�tƃ�	��/)�=.�>mh���*>L���wV>J�<e�����զ>�Z?26���h��==������
���b;��5>l�_>����m����>�W�����&���>��?5f����>��?�(�������>h�&?��=E��m�>uFw>�"|=3h@>�xE?��>?'?-�>f��=�w��.`o���>�B>��k>M
`?�8�<ѐ�]�z����j�%�ﳾ�ۦ>v�>,)R�Ó�>��=v�����{7?+>=�<�!
ͼ�]i���?{���V����=�:����>��>?=�T?��r�Q�����g>�[n?��=r�پ�޾�@A?2O�= �*t��`8�JA�>M�[?�Kp�8�M?����;��=	sB>)_?ع½#�����q?%X#?��4�Ēվ��>'��>"p=P��>vU���E��Cl=~]�>q��־'>:#-?D��>��>�S��f>2�hP��y�kk�>0�d�g��(��:8�?�%7�S�����*?�'�<��9�,�9P�>�Z�>U�;?��_��?�$�J��;��1�>,ń=(���W����G>�,����@:ʾ��?�>b<	?�+����>���?���>���	�n7!��B�>O�������~?8^�=�@fD�7���C�^YQ�ܐ�=��V��#���G����>U_��h꾗�߾�A%���=��x�ym���>K�UZ�>�)�2���	�={7<>!8�����b���0�p�=��W> r�Q�鼑@<>Xiv������h�dF�Ϣ>e?G<�B��H?��=8)����B�W>j��<ii3��}<��o>��Z?�짾���Ι�=)��>S��>�˂=d�Y?v&�=�w��D>�i_?�3������B8��EB�> ;?�4�(^~�Xپ����h�=��T>�2#=`%�>�,=�=���>��=���8}�j8=�‎?_�>�)�=.�o>��G�葌�	Z>D����P&;��=�+u*��<>3�I�FH>��<���6�2"�'��57��zN���f/?"M"?ɝt>|�;��'$=b�=���>�m3���=a�B;4�?��{�J ��y`?��ή>d<Ͼ��Ծ�F�> 7>T��{��#�'>���>�(G>+w��ξ���>�K��< >A�CT]���>�}k�q���U�d�x>�o�w�=ޕ�6�>�V�>_CG?�����̾���=k?nD��yy�O7>L{��]�7>p���'���I��=@?��E߾��t�U?}�?�@k:篹��w�>�<�>	-�
n��cľ��>�o�9�%>�N#��n\�直>#?�'Խ{7��CG�>ջ>��½< ��T�½A�>qV�l	�;ҽ�[8����&3= 	�=�k�>��b�@�{�q��>-@���׾��r�=^qs�ڶ>+��>%�&�+��K�:>Ѽ>@�꾢)���:�v]?�T5?h��=�Z�>&G(�k��}�	��C�l�?�?H饾�^�1�"��=��>g��>�&��C�%� �>Ú6?�qJ���9?�>�?й�=
H�4��>���>���>lZ��~~�I��=�S?�����>�骾���>{B$�B���Tg�� c�<!�=���>�ɾ <?�U?@y�=̀�=)�Q>�of��S>�js=�?��h>�B?u� ?��]?Z�4�즽�0�>Sw3?��>��̾ꜣ�}�?10���^1�-��Z(��Y����U�>h�X?�*�h/����>d��>�q!>X��*U�X�Q>�#�>7�!�A>E�`�V)9>�H��3žȑ+��T�>���>����}�����%n2>(�X�ܞվ/��=�
$?������=���=��>R���5]�=3_��7$>�[>Zk�>����.�>��2?��?������g&��_�>NA��C�|�����'V=3�E��s�=ks>�%>*57��ё�5��>���>&���ˠþr�`>��?��Ƚ?(<8��>Cg�ࢲ=d���]�=Q�;���>��C�;�)�l���y�>Z�A>�䑽 �V�3�>J��'y�ZBμa���}m�>�u�>3S��|Ʃ�Or>�!?��>L���[�?ĩ�>�7���(E���B�mP=7�'�u�$����>׳ >�N�i�Խ�h>���=\�]�w�#��?���>S	��9�.>�|>%�`=���<�f�>?����%�>sY� A��lg?�S������e�>�<'G�Q)?�o�?���eI$�f�^�ƅ4?�]���x=�#Ӿxr�=������=v�����>�� =Z?�~��ܔ�"l����J>E���M]��2�=��q�Ex7��Ԓ> ����\>�'��$�������� ���	���>F.�>�(���>Y���Uᗽx8b>�i~?�Z�=��8�iu.�@+�>��1?"T�<�Z{���>x>�(��Ѿ ��>��@��l}B�F��>5!%>_j&�ޕ$��SནKD?�&��_%̾��>��=u>�{?Fְ����逾�5?��?�P���:$h����>!�M��'�V�)���@��>�m=�a�=,5ƽ��=��\>�?��оj��>���>iB<?� ��M�s��v��k�Ƚ	���A�ig`?�?�,`>���7 P?�>l�>���>f�����=է�>˜޾(H>X�̾�C?ٰ�=9|�z����Hu��b�[Z�>���>�>�;��>}6�i:�g��>&2b���(K������L��2?�9ƽT8`>5C+����>�褾Q�>*��>��<�S�S��m>�W8?��>�9��i>=�=$���Z씾�i�=Ħ�>���=��S�#,ʽ/�<�Ȃ��g����<�.k?2�4?��>���>S�Y=3a?Մƽ'�)>�V?7�;�������>'֘�s9�>ف
>ʓ���i?���>�X��8/D�.�>���-=>2��)��Q����6?����^>uW>x{�>��ȾW�l�)���_>	���2,��F?�H�?͡?vKO������oKx?~1�<�]�{����N??(&>贕��V����>�+�>�4g>��>����ͪ<m���<�>�BS=|[!�S��>�`�>�E�=C��y�~a��#��̐��S��>��2?9���1��<���>�x�>7�=��.��QU�b�T=��>����ÿ>�w�qS�>�J6���x�a�!>Z���zG�W2�C�Z>H[��7�\=��>l�?&�(�_eU�*��� >#5����>�4򾵞�`��>c6��u��u��(�<{F)>4��=ĬȽK߱��>?4V��g߼~�ƾ�2	��;@�|�>������׾d��pC���b"��s��E>H��������ψ���?�]R>w#���.(�d��Rx>�B��(>���>���>Z�L������7>�C?�ڒ�w�̾��?p"�>�Խ��<�?>"�>%�;��(E���^P�=Jx>�˾�r
?O~�>�->�6�nPm�
��U>_)|>�����i��j�>����Ӿ�������G
?��=�"��Ue�	��> ��ܝ��֍���J?����9����Q> =A⌿p����w�=�Yk>V5>@��Z��bd/?0�1�X�༓־B>�-#�>ژ�>�=�⳽[<�����o?p'�(9��Ӿ�O>[��>퇤��h&��'�>�E�>�p(�1�5��<�r>$���@S������M"�>K'������PS��{�>�J�=�G}>����U�,?�$?݊�1L?���>Ǣ/�]��>u�??�?s��ˠ>�X���<!��?r�=�f�=]']��e�?9�ؾ����>=E��ut>
/��:��Mv�<�>v�>d�>&X���<Y���ݾFji>؅4���>q�b�M�U�!|T�4�ڻ&�x��s1�{<���)>���=	��YI	� 6>�E����=�$8�'���Y��S��u�v=2��>��S�^��_�H�FaI?��>�� >h���xRX��O�>�w�>�-�+Bs=�&�?n��>0+>�;4��8q=C3�<�;?y'��>��оb���@��=8���.>�e4> �?�⠿�������>�)>� C�&��=�����l�Q��\c�V���	>�ݿ�`H?�Do#��@?��G���S?���?�??ս{����wm?b�>b6a?����y�>ub?��&?.ڕ�ϣ�<�X>P�>59>����Ƌ4>.C?I�8??���zx�4o	?$�?=�zk<աd��	!�j�����۾�?�%�;�����@�N�����������=̜���b�7�'���=���>Kb���R�?4?���=�.d?/Q������������>�.?���=�~3�[c�n��>nlI?��2�(\⾜�A�p�p?�A?Z��>�>���?�w�>3?q>����V9�>F9��`�@�Ͼj��=\g}>����&3���?x]���;1.�>�ÿO�>��>��A:5�O����>t�G=iw	=Q�z�n7���y��=>+"
�`��<�ѩ�K۾����>#��<�hz��o�Te��*W�>瓐��Q���8=a�?Tެ=%�k^�8e ?ڼU��"��������>�^���R��u-��S�=8�+���j��󍾀�$?r#>�P��j���zƾ����>%-?d�տ[�b��/4?���~���s��>�GɾW��=�D>:.~��>>`X?���%��>�7��^����[>��>b�������>o>������\?Ծ.�/?*�Ǿ�'�����>�뢽�B�=E>�#u��_�>^M?�����~>DN�5��\>b��>�E��`_��c�>&�ӿ�]�>�?[Yu�H�?��<V�*=�X����>3b:>zө<s@��Mj��K�>�M�`�'I�>�g?�]?>��<鼘?Ud`��mb>��T>��8��m��+[��Ց��+��o��>�������>F��>�a�> #@�V{?�'��H~>��X�>��?�N�=���8#3=���=vi�>���>áK>S`?j��?W�<���R'?�N~?��K��Z������'�҂��o�E���a���н}�9�}s������e�6�>�-?E��g��f?Ӹ>,]{>�/0����>	�Z>���>���{�r=(��>�r��gU��Q�>k�Ƚ$b���䠾,I�s�ƽ�J=����b)��9I>R�{?Ded�Q�=�U�=�`˾e�ݽCL|�ڃ}?__��D�=B�n���w�?�;���&?��k>��<�aj��]�>]��>�,h?����v�>�p�>؂����?S ���<=Qf>0j�>3���Sǯ<��쾨�o>M>���ݾ�/�����?��!�n;���>�L8�����'D��>�6ӿ��>�6w>�hk��L�u�o=_� >BM�=�L˾Gd(�Y���?X���ʻ�2�=�-=�����>�f�7>��%>v�/��E���/?��ƿHf ?&��=C�½a��>�c���ON�7q=�?F�=@Ÿ��z�r�>��>�<?��y>@�>�����}N�!f���ھH�S?�=�P[�z�?�'?��H?Se=,!)>�.c?�ޯ?Nn>YqO�:B>߂�?�p�=�[:�7�ɽ?Q9?�θ=PW>7���D;?�A�>��>��A��$?w�s����=3�Z��Ce�{��>�%S��B?&ե�Dn�= KB>��?e�>}m>���>J?NO�?���>hQ�<N��;	��>��>G�/��GN>w$P?H�2>.�H?c.J�R ƾA^���`�?�Ԩ���3��Ӄ_��!���QT?����k��G��>_��>�.�>xA�=��=	W?q�P?�s>���|��>�5��7�=8��>'8��/���Y�M?>��=8wB��6�c]>ʇ	>0��<F�O�4=���>��=�u>�O>���=JW���5>�/�"[4?������཈L���?XE>�mF?Q��6���Q;"�=����-�Ӵ/� 7->�	��
>���ɮ��b�;G"��Ġ�>]/>
��>z����'=�� ?t�>	*�7,�>c_�>�鞾k�b?{���N�=U������k���1��U�+��>4N[��I�S\>^=�?0DZ�u$����s�*�B_��mu:�2�?�Oi����=� R��ߒ��e����?���>���<�Td�E/Z��鸽V��>�߿�s���3����=}\��[��>SG�=���>���L����0?�k,?�󽿤��>�&���R��-1��,���(�>M/T�@��>w�����=�о�D��]���%2/��辎�D>=�D?4־T�/���>�k�>�;]�q�ҾmZ�1?�&�?���J�� 6�?��غ:�����u��nK���:=��
�a��g�?֯n��c�#J??�Y�
7��<?'������r�L�����?2A'?�dk>��9?�U�>��>�����?XĽɞ=��K�^�E?��r=cL=m�>���>أ	?�l������)��?4V>�hF�@˫���=�8��U���#���K=�b�>sY%����t��>�8�=��k?�/���=/н#�2?��/��=}up�z�׽�@	>s�?t�/��	��_b���>���q$=.!$?za��� a?j�>�� ���6>p�:=��ļ13�>��-̾b4=9�=��B�����Kq?Y�i>2]�����R(Y?�U�>�3>�o�x@?� _? ��>Xe����>�p���h�>�&����?�T�(��<��?��Z>(z�h*?��������X[>�W�=� �����"S��%���m<?�C ?�O�ۓ�?�?�=RF�����}W�?�n����ս�X����>���=�@d>KC*��T?v�Q?}q+>n2��۫?���>�D �w����>�Q<��;>����M�=��>ɤ�<�>��D��?fޝ?RþS�?�=>V�
�_$ ?֍>�o=x�>��>G�۾f$Y>�?bN�=,�>�>(?x�J�0�I�
��=��.��>��>�ы��Ѿj(�3aپ�
����+>�d(�S"�c[��qG���>.��?���i=���~��>*�?o`�>}�<�㡩�L�?=�?��D� ���y�]<A?d�?��>�)�}ԗ=@��=S��>��L?5A���=\ı>���>1����Z��i���ƾ�,W=�%�#<<?��Ƚ�N���#���&>�??W��z�R��4?��R?�8>K�����?�4K�Pؘ>|�+��Љ��\?�7忕�\�"�5=�	�=7rE��J�ҵ�;�򒽇��>0󓾘'�=�{>W矾�
�>�#Z��X�V&�>���C\�������TL�j�Q��a��VU�zƽ2bq>����il��f��b���Zk�Y�>|�Ϳ
�!��y׾_b%�Ⱀ=I;*�	�׻�z�>�\>����??�>>��=�a�վpϾ�� ?����ȡ\>B7��%��>5�]�T��>��`>Y0�>~X>��}�<���>@�8>�׾7�K�H �>���>���O���?�v<���=	�Ծ�`i?�U?�B>VB(���W���>Ơn>��>�_,���`;�ѕ>�f?�����G]��L���c�j�+����RO��*�>��L����މ�bL�>��������>��"�J4�J5�=ټ�㾉�R�g��]���5�c��>����M񀾥So�@+�z3g;R��"�?lO��>'����)?��'>ʪ8��o�>ZW>����|b�r�ž�J���	@E�W>�Y���O-�f>���=@����+1�e->�ߝ>N��&�,�ܢ>.G�>���=��=޴=
�C?A2�.1+?ёZ?��>�m�>�?2p;�?�#�>_i�=�@>rC	?����4�=m)u>'�>��2v�>_5�><�/?���:����<6��?�2���a�޾A?���;����&��R=���,&K��1�>4�k�/4�3w]�'����λ>������藾2@�>4+M�A$���>�5����˾���>3p�F<�]�םJ>Ľ1>�?�̽��پ��x�f'\?�.7?��?sX����1?�c�>gis��磽-�
��<�3�>=J=�z�о���Ω>0c�>@�+��a��d��?��j=�2�B�p�
�|=�x�>���=��ؽ�p���hu>jc-���p���3�>[�\���	�l>�;.c >&Q�>gTc=e�3>-[�=^�����r>�nE>Q��N8>��W=�J9��ڠ>��O>�a=\�ͽ�9���;*��<>���=�9˽�Θ>J� ?SW�+^Խ�s���>������S�Ͼux�̖�R�0>G
2�q�<�&>�)<S�)=zv��K(<�m�=0X��i-�}�u=��6>�:��t����>o\���ڽ�!q=lA�=�"J<�ݣ=��=� ?ܡ��C=Q�H���g��>��%�ٻ���>��?�]3="7�=�/#><X ?��ӽk�=Ձ�����>bjq<�����`�Ա>��9؋l={���co�>\���-+��]t�=rr�溜=M̲>kh�>[hK�DC;����=y�_>������������g��L�`E�>�׫�)���W��1�>�^併2/�����}�=a��5������>�b>��J�hϚ=��%?�
���ԯ����9�+>5Rۼ.)�������>�_s�!#����<�v�>A��=�퟾�W�<��!=�.��MQ=��^��/ɾ�r[= �>@>��Θ >��;�9+>$M�@6��,���<^��k����>��վ�x\�`N���5u>c��=�I���_G���C>�$;pJ>���'����>?(Y�uK��[W�=C-�Q��<���w��_=��=Ig1>��=<̮��m"<�?N<-սP ��;WL��/�����7o>I3��Q|�=ѷ�>� >�Q<Q½�}㼟�&>�]ҽ����"<�$7>bͼG�ͽ���>k��>>]f>�:�=Dm?S猾Ay(�=t!>��=1�>�彆�⽪_��'N>7`�{;.���0>Δ�>(7f=[��=��>qػ�L�\JX�{B.<��>>�Zڽgv4��E>m��>��>M��=��>�����"ҽ���=�ܽΕ3>�}>��C��������	�����2k�� �	B���I�2쭽H�&�`�I>�=qcK=�o�o�<��M> ��>����=}�=U .>'q���*b>��>��=�g��k�/��<�L>M(>��1=��%�Wg?�Ğ�5b���<<��=N�y<�L���Е>[��>�ٽ��a�nS%�cD���Q>��5>Lٚ>����>>.�>�d�=2�Ⱦ�9�;A���⏾�`^�E�l>������>yC�>�Y¾2p]��@�|N�>��l�E� ��t����>	>z��>��>6��>�7���Ͻ)�\�Nz��dz���(>[�=�\ʾ\���"�<��>>��P|�_%��I��=Ⱦ|T�����=�-���ʾk�v��O�<@,>���xk�7�,>WO�=���\�ƽf��#���P ?>� ���=�ܛ>I����v)�&:��][ >�P�=RP��fOu��a�>��>�T?A�->z�>6-�@�^�er���gоGץ<�� <��E���L���=�#D>�y">����r���,l>.BC=�v��+����>S!;>���=)������=�#p>�
i���h>LsT>3�W>M,�^^>$��>��/<��	=��>�������>{½ֺ�����>���<,��=�Pl=<>��:>�H�>���=�"S>��M��Eh=�2�>��>�'>]��>y]=�*�>��1�v���@����S��E�\<�H�aA=��>�����}�>���=!�<���)�����,>c��=��uNR>�	�>���=�b���>� �>�7�a>�>������:�H��>���<�a��	nz��1>�/{�w9@��f��I�\>��<��&|�>Xo4����5_��������>/�>ΨE>�渾W�z>���=�o�=vӶ�$y�3��'+��Π���ɥD=W�9���^���9=7��o�^͵�t��<_c>'����?����=WQl>牘�	�)>�'[�<%n>��j>T����ϑ������h�>L:���ռ���ڑ>m�<J��=W=EX�=��T��5)��s�K����>-�;��漻yݾ�����?����W=����@^>���O>��������I�>fIT�~p��OP�|wW=Vǽ�k��Rӽٵ��н>�-�	�1�`:ս�}>	p��g�(�}�%���8=UO�<� ����T=���=�����9�=-ޖ��o���*��r����!�����R??��+&G�; �B��=ɀнy��|�ѯ�>6��k��/�'V�>�K�)w��J �O��ƕI��#e;�\��i�)>�>�=�=��ӽK�[���ؽ4�|� ��,c��׶�B����p?bϮ>�Ay>'d ?���݄N��,'�x��>iv�YE8��=�O�>��X>j>Qk�5 f>�)c>H���T�=�;�>27q>��=}ý��6<�>.
۽�(����<w�,>m&<�-<�ނ>��s��:�#��>_>�ܾ��T>�&P>�/=_��M�y�	>:*=7>K���ྜ�A<��_��N�=0��=:�ļ������> >��
�]&%��H�>�ݰ=��?�z�.��l=�g��/���5ʽݻ��XT>lp!=�|�=rY���Ϲ�)g�=�w�>�#Ѿ�->2pe>��H>���K�0>'޸>yؐ<k��7��<NI���G!>�Ds>�	��|G��)s��c�6�$u>j�F�z�ڼ&�(��p�<�F��lM>��=(]>3�>E�<�/�ha_��!t>�p�.i��T���>is>T>�=R.X>��	>26�=�'�s~�=�>�j̽�s�����=�k�=I�B�����>�Q�>��z>�7�>��>��>�L�=-���Ͱ>��+�{��=��>�XH�|��>	�=u�M=J�E=���x콟�Ͼ�z��<�>�½�����<��>n,z=/��V��=L��68��+��xW���q�[O#�k8��ׇ�ޚO>*��=uvz>M��F�<�-�>�?������'����=���>䵽�<�=���=��>W�2�}AA�eϮ=��O=����>�>����b9��D��<�s�=����k��s%����8޽&꙾�1�>S��=|�$<5z�)���K�L>�d�=�b�2��>D��>V��=��'���>;�>Sd)��ݾ��=���\������v]e����=�F(=�\���8 >3�%><Ὢ�h�w�e�O�J>����d�q>c�������K=�Ru>���<Z�꽪y��C�=���~{r��Ј�Ǭ>_'U�i��|�>�mp�ߏ�=��ӽ#B~�VI�=<����*���
���G�ـ�>O�x���~�ɜ\=]W|>ϑ���a��Q>���wfk��0��Ⴝ�,�=���m���A��=a�:>���r��Ni<�.>�ӱ��Ҿ�1>�f=J�=�˾u�D���j>��7>PF����B>��>�y=Eѻ�`Mk�hv#>iP�uyv>�6��
$�k7�<�a6><�j=I�<��:����=qM������Q��y�=��A��!1>�]>��&�X�8ƃ=�1>z�=>��������>��&�������.�k�+>�#c�c�ھD&X=��l���<E��Q=���o�����~��>D)-�.�Ƚ{ �\!�>�0��>]�w>��%>�9�>ߙ���`����Ϻ��>�ŗ<c�a��y� ��>�[���<ݾ�0��
�>�jl��fa�4o9>�{?�d�=	�<��1?W?9�@�%<��>c�+���> �>�Ǡ=��=~�>>���<�?��A�=���>k}S>Wa0����P>�;=]]���4���\?�����=�!�D����>Jμ��,���"1�SH�>ơ��^��6u����~>�_>M�����^��X�>�k{�����W����>����`J=�-,�^����c��6r>��n=� ��PN����=�n�=o��ۯ����>4uj�㭟=��������z!>�'�<�4�=_�FC���<[=�Ia>t�������/�5�>�����=��[����<�n/���?�-7�x@�>�pG?,鉾�=���l�>�BP������ �a%���L="�t�7�-��v?J�?N[�?�x�>M�=��>��@�	&?GM�<c3>�
�=1�8=���>��R?F�?O�x?� ?�:/?�PO�Xf � ��>�I����?R�?��1?|M�>ML��U�Al9�y?�g+�UFV>�h?�@D?g�>s��=´��dܾ�M�=�2^?��"�B��T�����3��Y���,>�a�=�Ý�g8����2�n����'�^�?��?��`?�J�,�r������?���jؗ>_8/���_>�u0?�/�?��"?F��>m����>?��>���>�^��c7߾��
?k��>�ڽ(�\�d����>��?�o<��Ͻ>����L�F�|>�q.?�v3?�9W?�:?5$����t��J�=�ɐ�\�>Hc'��"��s= ���D��$?}&���mA�����ٔ3�2�=�BP��ϒ>}���N?�ܵ>���u��>�Q:=����}��>^�"?�� �#���_���I����IH����=[��>�D�e	�����|Z�UL��-����?o=IL��A����zR�>k ��V���O�w��=m����=g�����?o����=���=Bj_?���q��������>+Ƀ��
���r�2ɽb邿��۾��(����=宬�=���C�hc?C�?��V?���;�݅��S�#<J�����&߾�K>5f�ƫ >x)?T_(>�(?C,>Bx�;!�I���>��̼��l尾G,� f�>'�>(�=>��=GR�>8|W?���>GyK?�K�>������=���=�F{��	��B����?���<h�߸�����N�U�v����>��s?	�,?i��5�G��>��Ȼ�G
�<�a=?2�_?�_?�ӱ>5Z���>�wA?��$?�Q���>��>�>i$�>��>zE�>�mr�.��x�<�
��bJ?����F���O;�=,(��(��=f��#����/��e=w
f? m;�?P߮��ѹ��q����>�Q@?��[?�A����WJw��K���.�����`�L��q�>	?��-�����j�dz�����ӈ=�|>�쭽S�H?鹗��j?8 �zK>LД�Q@?����/~)?CT?����6]þ�>1M��8��7M��ݽz�)��L�>���>j��<J�!>�����=����u�>tu?�G?�m9>`�>1�>'�>�zq?��=^�->V�⾬h >�:V��̸>Zľ*�a��s6?ǑϾ�O�����b@�>8?�?�_�=<��>����D_�\87��žl�?��Q?:�=>���M-��L�0�yO��>�����N���Y���C��<�Z �%�W�kh�>IO�>	�ټ�����V�>9X���߼}�>���>�6?�.�>#�u>�#?���:����ջ�^����z�1�>{��^l�=~K���>?�*���V���>c�>W�?�%�>ɚ?І���>��/��T��U�?<=?���>�Bξ��[>e�*?���>��s�~,�\�&?�h�8��>*�׾���q�ľ*���Ծ�ey���?,}�>��? ~۽iZ�A7�v�?�?2�c?k��>��f�Wm>:
�k^�����>�2�>k��?+�>;$���j��צ�<���,�K��?���>]��<}��=K>��';�V?	�?-e�=�8/���"?ť�?��X?w�+��K��#�?��8�A�?��>*��>���>���>�fo������3�>�>ss���/���#����>[�>�!��̦?�r=>�q���5�(i*���ݾ���>��>,jW>z�?��g��v��g��bM?x�ȼ�u�>��?�&)�����u���Jоe[=�}��˾-���L>�[6?H3�>��}��5��@�>��>F�:=�J#�b;��S�?x\6?����0��y�	�&Z=��/\����=NC�>�5>�z���#O��i����?:��	�q�L��14��)_|<o
޾������ޏ?�hB��.H�7j־q��>R��?^)�?�̾��ݧ��:��O��ï ?���g���!��g�>L_
?���Pھ]�<�o.?�g��_�L��vh>�MG��ʽ�EX����V��{敾�'�$��=�q�U��>fhe>b��?�lؿ�U��o��z?ʃ�>��>��O�� ?��/��(��SX�Y�?�{��$V�� S��B�m?�b-��"��<�l�� :��My���؛��Q�uu�>�H?J@>�{%��e+<��k�V�����O��~����=_b0��x*?7pl>>S�?։y>
�~<�v�=/&Q�赂?�A��`��&EP���?١	�Q�l3r=�i?�����`_?-��+�<?'�n�+�;�����*>0+=+���@��d�ǡ��=�>Q�;��諾ύ���u�?H �Y�>��0���>}J?��"��-X;�w��7.?�U�f*��R��x���`B�>9?|탾��@<Yٟ�����O?�L>
\v?�Õ?q�^>��f>]�|����>�81�zЪ?�� ?�'=����H���C
r�32�	?k�Z>���>�qC���>%��>`.t?T�!��?)?��>?���t��-s�������@��@���"�=@?�`G?k���ڽT,��`����T��V�G=@>����0��W�^�?���?���>jƴ=#9]��A�>�o��ڀ���^>��?XQ>E���*f�_�?B·�>��=Ƚ��K?L�xґ>�c�-ľ�i<������>@�:?;��>$4��p!�}�=�J��>�Z>�.?�m?v#[?v�?�i�=�R�=`'�=�J�>ݛ=�;?�A�>T����@=��		����`��Hk�Ձ˿�3��m?�>����>-����Q��9s�um>V�b� ?h�������������1���n�td&?��:?v	<?|�!�f��cL����?��5�`t�>�k�>i���fK� ��?Z0���>�8S?8��>�|\?3����B?�	%�� ��<L?��*��f2?��`>P�?�+����zjH>��;�T��l�>V��>���u�� s8?F|�?�N�?��$=>�?�GZ�̸������վ{ ����z�����;�=N�>`�<��6?�I>������ɾ��*>i��=k�#���97-?��>y�=��>������}����>�>�>䨿��;�d��>'t>*�V���>9�:M`�s��b��������&��~پՅ�'�<;㹷=�vq��!���~����?w"�>L�L>H�y�����<!�j3�<���>���@!�����|e>�YJ?�ǁ?L�?> :;]�ýs6 ��28��86?ɢ�>0H�=����������>�
?ukE?�Q�
�>1Ŀ>ߵ+>�M�žV>��f?i?j3M>j�?�	:��2����M>q*������X=+�>�<"��ſ����м>!`����	b>����H�"?�{���g>v�*>`��q,�������>#(޾���0&E�w|�>�>�凿]��>��W�Q�½����?�$=\褾oŖ���>r�^�����M,�=K��?�����?B4�>�@?�*?�@�� ,>�B>iA3>�1������nZ�%s=*ֽq�I�c/��SE?r�]�����>+�Z?g�x?���>PU�>�F�?]���H8>0~�>�$=��m>w��>ʍ>?sN?���%*���Y?��D?��-?Lz?k-�=��m>���>8Q�>I��>׎f?�b���:d��짿y6?���m���N>�&#��>����(�=��;?������q������>�`
��ˬ���7���?�K'G>�!��۾{���O>���ϮT�'������G�!ʚ=�,?��>��>��˿Vd὿�g��f"@k̚?1��*� ��8��j��Ⱥ=��<~S?���<�9�>�>U�'�s�o?F\C?�rW����M?>����Y_?����-?F+�[����-�|2��B=��j�����]��F<�=N�g����j`�H��	��:�?f�>t��>�ſ>�9?��>	�?k�?��&:����	�>y��?	}3?Xbm?�n�>��>��>x
~�4��ҵ>�*?��d?Z���ľgQ���ZJ�ڌ:��ڮ� ��,��m�>U���X�?-�?g�;"����o~���%�93�;ʨ�<;H���=�K�>�+�j_���Ow>>о���>���>�D?��&�:m½1>�D�=�4'�K���iE�ZnD>^�=��W�/��_��̢?ݞ�>81?��>��O>�$=>�S�㕐>�*i=
@�>-��Rn?��>Hh󾐅 �$�@?Ѡ�=���>>�8>�C����Ҿz!�>��?r9!?���*��>3�uv�k��[D��Td=�3�]? 8þ%W��Ω>#�C>�%9>s鞿/�	�L����$���H>�����?��>_?�v�>��>-�3��Ǒ���۾�D=�·:G�#�
�=3>���L�=Ղh�oy�>l���)�%�3��󕾉�N>k�����o! �ԫѻN�>�����_=�='��~=(��>��N�`׻>;�O�v��Uzs>e"��m>)���>Bm������Q��A��}dl�$V���ɑ�k��>ƴ�A�?�W��V�*�Edp>Un����=������>K�U?U�W>�3�<�N.�xTw�^ϵ�M�����=g�=2�ξ!V�>9l����?��>�O.>������"����<d�=���>]�h��>�v>��9>�=p>���?YN�>K��>��>�� ?i��D�I=�44���Ӿ�O������o��cV>̬#?�^�?��C܄���e>�f��엽X�x?R��>�7N��i���������h>�K�>���?r�d?�?/I��F?Lܤ<��J�5ݳ>��Ͼ���K\���Z��k��>�,�l-�>>}m�)BB��Xg��a����>��nHj�T��>�&��x�>P�(�~��>��?��>�n�=��k=_$?���½5����d>�I���>9>�� ��DW�XZ��QT��X$��RǬ�{�(��>��M=����$�ѾP��{����=S:����D���K>���?�t�>ꆈ�6��M��>�y>�Z���2�=3���?�$��N��J�K=��?��˾��>nD������?�5��Ș>�9B��fu�6U���҂>*������u`9?�¾��fH�=�Ծ&�'�sR��X����M�~�g?䠿>�v������ŷ=�s9>_���[������\�>ϵ#���.�`?�+彗+O�'��x�>���?��=$/�=NE!�3��>�����$����>�6u=�#�X_>�����)=�7?��>xbV��ˁ�[- �<�?��J>�>�>id�?Pa?R\G?�.=�TB?�;��<�>ڂý5��=��8?rw"���!?��=�y.?�q�>d��>��<��~���	?I�J>�k]?~T޾�C ��@�z�z?���I�?>�P?,�����^��=ɵs>�޺>�,=��=�����>����|b��17��~��<,�3>�`�>��)?�ۻ?��?.B?t��>�)�n�=�J<�܇?�=�%�_>5j?�+?��>�f<�=��_�?�\u��Z?�ǉ���C�'�Ѿ����H�>��V�L��\߾�Z�=�X��h?>��=��>Z~>C$3�<l������f5?H��>��u�WG�>O_c��<��>��r�X>��N��$>Z�r#���<>�w�>��>'r¾$Z���2S=lv�>yǜ>�6?z�D�[��>�D)��P���8�>��<Sc�?�m"?�&q<L����05�3���w��Z��>,�?��������T��9&��¾&�o=�,(>�J�=̚��� >ղ>���>��������>'��>i���=���5>��p?��n��5Ƚ�Ŗ��t>�����>��s>���>�N��g������3�>f�׾[���}����M�f� >m��=_j�>A)���>/Jt����c�Ҿ#�c�T�.>Q�n?�'�P����m�Y4�Ζ�;L��ޞ>s�>N����`���e?�!⾭{v���-?�z�>j���'��>���=�[�`�>��>��?=q?��u�\Y6�A�d�r7�ulU=Y��2y?b2k�gn�>�XR?�W�����9��bI?��)>nSǾ�k��z>4�?W�>��d>��k>�	q��a��}�>�R�J�1�����~\t�0�>�Қ�=��>��|�Mw�3WھR �����S���������7&��\�>��ɻ�o�>��,?�ps=tJ<��n���>��s>o���z_ �w�?:�>��G>����V?js!?0J>�,?�F�>�s;>�iľ �a�&H�=8Gd=�4��#\��_�=B��<�^����6>C��>U�"?V4l?��?���B��Fb��e���R?�R�M�='9���?q� ����޾�Ar���J>���>�?>Z���,?�^�<
_�>�;>�� >���>�3�]��뿰����V���{������Y>��O?{i�?�;�=�^?�+�>�6*>d`���	��|�>�v>�ڽb�c?�4(����>���>��>B7?�ܰ>����Da�=�2þ;":?j;��p=�G(�h���
��\�We���7��>J��M�j>�~E?�u�>��ھׂ���=}�>lVY>��x=�{?�q�>�v?q5��0?��>����Z����;��+?��t�Ѿ�H�v��>� �>�,�>�bS?Z|f?Ue�>�襾-�?P�->���>͈|���I?���>2<r?fƎ>Ԝ���0?RA?���?-�x>�G?=�	?��<,e?�?�<���>����QT���X=�Zr>M:?�L����m=;�%�u�E����>G9O���*=Qk���%�]�����=T�Z>_�Y?�IV��"$���K?�dH=JL�nY��c��I�e>�@>��C�܍\��gb=�p?��>W��?�(�>��*=�_3?Y�ƪ�?4ľn|�<�4����.j�=Rk��}������@�>�q=�^#>V�?C�=���>�5=>q]��l��Q�Z�H�:?#4�>�3a>�,�=���q�J�C���?��0�m�P�ߢ��״�>u�>��=i��}����� =�E�ل8�ް����M>j1O�W?ڦ&>&�>�G���xW���<�0)վ}��>3bj>��?>'46�q�f�����h4��O�="2m��K�C��E��cC���нC��VAJ>z�=���=tgt������K5��7"?T�0=��TG��=�>�4��r��! �>U>�9�
��߁ý�
�>ps?Sͩ�H��k"9;��P>�Ȱ����=ќ�>i`�?ʷ�>�'����x?]�#?E�=��;>�t�v>b�꾽���x��>uy> ��>�ڙ<=Ga��=/�P'ƾ����Ӵ��S�=N��>��>�($�V����7��l>#�|/>��@�>�?U�=O�>ohc�?�X��U�Uׂ��4�>�ܽ��A��;���s�g��<���:��=ץ��|�>b�u�\,j��-?M��'s5>��.����>�X�[�x=�؛�Ռ��y�2?k���$�Ͼ^���'��>�Uþ9�žE��=��e>�Ӿ�&���Ҿ>K?+H�=�t>�1<�K�>O��>�޾J�?�S;?��Z>\z�>>��>䂖��䴼��=@g={\�>?K����?�����v?�JC��BL�Ҥ[>9�>S�Ë>����R�<��Y�M)�>��%�W��>d��=U����y#>[����EM�W[��3C���"?E�Q��	>)@Ŀ�����G�&��>�����;>z�@�\�A���;?�@����>?<��,�P���PR;��'�>S�(=d�W�˶�>�Z�>�I.?q!^�h��»t���]�Ç=>���?+�>A�P>E��#���9�r?�Gg���Z>ޛ������A􀿦�4���{>D�zQ?�H����`=���!�>�*�=noZ>�rN>�2>��,=-�=���e*>��Ľhh���qʾD�{>��۽���H��ªU>eߎ=O�νõ�>�>�I뾧@!>�?�'�=8�^���g>b����F���T>�?=|��������d[=��9>.��<q�2�N��=��>��<k<d�Z=��=3F�*�}�؄̽����l�mt5>,ʎ<��W=�'�>SD=������=���<<�2=�)ۼ�"�����f�}>ߡ�=Z��<�j>d�)>���=+^6�Ђ�>�&X���	�=�P�>2>J���v����=�Z>G�I=)��=�s=���>�U%>]�b�=W%?7e㽐���> љ>�:��KսBI�<���=�(H=%��=�x��*2D>Uc��Q�=@X�>�<��}g�G�E>���>����%��*&]=��)=^T���3�ˢ�$U���/�4�=�_������~�1�>rtC�����@Ҿ���>�>鑰�k˘��΄>�ӎ>�
x=8����>0bH�+�<���z�>R ��N��������>FH@>)��8�I����>X?>ի���伅�Ԫn��I>�l�2��=�*>�;�=u�	���(=��>�H'�� ��޽����M��$=}��>ꥑ�*�>��<Ъ{>����I�1&澞'�>M�<蟷����P">')��dt="�*=CSԽ6��=�y���r��ndr<@.K>�8>�b���c��I�;�|��n�Q�V����+��ϋ��Z>=�w�~��=�->n��=�]�����=���=!�)�k�ý?�<?(F>b0>U0=8�8>��=b!=���=Ѕ�>jd	��19��J>�/���.�<���<���M�
��>��{[O���J>0�c>�?=�y��y��>0$$>�9�&Ng��m�� >�9�<����1R=�xV>+<>��*>lU�>�{�Դ�=��=F���ꪽ��=�l7�����->d4��E����������c�<ܽ_�:z��j9�>�c��X�=�v���G@��Q�=��?�4�����֌>�F�>�9g���z=P�v:�e���>��=M���6����J.�6X��:��� b>H@���9�fM�"�w>�����=�{>�U�>�w����<;��=4u��ah�=i8>��>����>qq>����vĊ���y<����!����l}���0>D�3�������>�d4��Ug�&�����>�Q9����;�.;�2�>C�Z��]�h[�>���>k�N��}Y�;*l=�9:�P���hU>A�\>Cp�Tg���� >�}>q$����N���;�$ʊ�c�ʽ~���+=�I=�Z6���6����=	�}>/��<Ʊ&�!����\>���;}�n�����W�mܰ�F�>J�$��W �:!�>�+>c"��`����>9�!>j��<�:���n_=yN>c��=�y{>��>F(��y/-����Of�yx�=��:J=��e>F��=x��>7�}>i�=bj�IL-=��>pG��ľ=��>�풽(3�:�-��m��=@��=X�?�ܮ��J"�!ɶ>�s ?ֆ����=Q��<of���AG��~�<�M��cS��0�R>�TӽB9� �7?�8�=��=���>�
>˞Ž�,H>�`�=���f>I�x=�	�=ޟ�)��$u=t�ͼ;ʠ>���IQ��zY��g�H��<��>�=�<�M
>����b�>@ ��\�!�~�����=FR'>ʪ�=_]�ÍH=��>*>�%��)$����=�� �/z�>�#����=4��=�>�W/�	Ӂ��ߏ�]�N>�y�x��pE���1>Mo�=\;�=m72>�� ��=���=!J���">U�>�o�>�=�"�=ӛ�=�2ٽ�Ǝ�hO{���=�����х�)�*����$�� �龚��=�`>PJ��f���HZ<�##>�c�=�
$=�L*����=�˽.�5=}�%�o,=;+>��Z=\*@��1վW�>V�9�k
���D>��>�7��iY���JJ>�� >P=?���t�sy	����%50>��5>V�ԼmT]�q�5>bj�=������T=yz�=w$+>#���0ʽ��"==�/=e�5�>=+�C>(ew�9{n���<Z�=�H,��^���^���m���6=y5��Q(�=T|=\�u>�.�>��"�<{>�ZK��	U������}��|����\>F˽ڻ�`C��i�>0^$����>�����>�n�=:�o�o����>;��=yd��ѐw���5>ْX�j���V�<H�m�y��?>w=����f��G���>]a��P>�������l�Q�}I ��	>�cL2�ڷ$��Aw>�I>�� =@�>�����Y+����M>���~k߽�u@����=�M�=�d,=ko�<��1>tď>�u�=_uL=9;I>��=�C�]'�Em~=��z=�A�R�+���޹�t>�I=�P+<�,>9�n���=�ϝ>�iD>�~���<�Z���[��X�� ,��"B�g������H/���H뽲�G=��=U�s>1�>��žδ�>f1v>����sZ{��Ep>�=�f���k��_#�nd�������	��+��_N�=�#"��5�=$?�����q�=M+?N.���Bw�>�ަ>6|����R;��>�ذ������ ���=�����
0��v�=ͱ=�~*�5�K=3��z�;h�{��2-���l��l�;�<�O2>O7=���<���>SO����ʾ��S>d��e�ս�Q�>YG�=xw,>��S>5I#>�n>+䅽�����->2\(>�ؽ�
�����=^�򽖏�k`�=tI�>8|�=q"�>xu}>��m�������-l?꫼������~*?"�G�f�=���=�(��'���&Y>p�@�+"r��S5�L�>P��>_��>�����v
�*c�>ʐ=�x����r=�-�=Zپ��s�k|=�5(����n_s=��=�/�=̒+��`�>b��!���/>��(?~y��Ô+��w>��>�6��8�>�|>%$V>�&��,/*=���=���<.d(��^->�>�(��׍=��>J̘=<�R�-|�<�sy�ÀV��`%�g�� �x<+[��A+��鑾5�2>l�>���=x�Y����=�ߕ>���=�5T�F���S<?��p��|�<dK��[��ЫԽ���=yh[>;Nv��d��^W�<�k=���9*��?KF�@���a�	@�>T=�<J�=hQ>�o>�����T���bQq>�$��a��?��K�s>3;���h�e��=lI �iS�=)��$����=���ފ���\~�mS�<������"<��>�F���C��j�=�$�cɋ������|�>���A�/�=ɪ�=U��'(�=S��=ǆT=G��<�_��z��eĘ�>?�%�ƾ7E>e�����j=�3��{�=!�>x�>��ʾ����鷷>b3>}A���'N������͚��>Q�[�<��:>�W>���.����0�j>K����N��bݷ�L�M>��Q=[^�9�k0>AJ�>BG;��P>طe>�*>�ܱ�GZ\�Q�6���->l��v艾m�;��>bΌ���۽ȝ=@#:> �=6���:��>����Ve��T�ֽ�\@?�nA��z�?:O>6�>2'=I�M>���>�`=�Υ>�����i<�����>�������;�D��>.FZ�T]������dV>
P=>k">�c�=��>��!�����2*?/+��8�N=���>�����.<�>d�X=�������>*6���<���l=�>_�F>:��>8E>�M�>��3>G�=���6��>��+>�����^RG>�bE�'�z��~���>!��<U�u>�Z���]�>�>�=@����%���>�@=+Ҩ�3�;[ۖ>�h@�V�ν�pI�l=C��O����<rᾊ��=�P=`G���0�;���>�pG>F��<Y%���k>�Q�>�[j>!.�O�)=[π��������>�H��	6��n�=ge?S鵾MA���z�>c�> Ǿ�pm�2�Y=]��=��>'Xc>�z/�"Ͻ���=s�U��=/��#��HR>�뾮�m=2����(?� a����Xɾ�Av>N�v=,�)�!d�>_�>�S>j�4��>??�=��?4�<?$1�2��>����%�%?Z��>0��=ɢ9>�j.>Y�+>���=Yq�=��>cV<?b����>-+2�y?>��0�0��k;�-���#Wf>�	=?,E��u��>��=��˿�=��=E�|>�&��bC>I��Ҽ�>0k�:tY��`=��U� ȼ�"w>
C>8�žfSH=�?`R�>�(����`Q'�?�?��վR<a�������B���>�R?��=�_
?y�_=���=��<>a�>Q��>t���H?%AF�� �>��R�>j/����>�E�/�|=R��>�T��2�:>da�><�$?j�??��|�>���م>*4�uN����M4�[,#=�LŽy8(�W)r�23?N��>��Ҿ5WA�Δ�=Ǉ��=���q+�>��d?+K�>�q�>U"k��$�=Tm*�`R�;*��>��=�|w�3�3��=f:�>.�E�<�vi>�S�>��?OE�	YǾ�9����=�q����<9k<�ް?�&�P ?�?�t\�HN,�k��^?��kٽ*
�<�s1>�/�=j1I�>�q��>�7����6��i��"�4�����|@>K����-?�̑=j`���U���Vi<���(�=�ՠ�q���A>G�9?���>+����>UB��n���R��N�Z���o>3� ��#t=	M�>.��酬>d%��Ƚ|�/���B>8J�>:���c��|P}��>���=���$o>yѢ>�w?]��<�3=?>^��d>�=tݢ��r�<^��������ݽ@��>�Ѻ���L��>���;mp%>�I"<j��>�+>�#����߾*5q�#��>�C�N�þ4�>�Z�>�S�>�Q>��>���=���>��>h�^�B�M>@;q>�� �>Z�w�;E*�����E�˽������>�rӾ/�����-�e�9L^<��
>�Aʾ���=���D	5?[T	�	6?X��=�Vg>1ޥ�$���?>W/�;_�ƾy����x>Fٗ��Ve��7k>c3��x�>U&�<�g<6�:����>�?h�'�#�[q�>��FF.?�� >٫�=S<���R>���hW�>oȾ= ��]d�?_�>�tɾ�D@>S%B�j'�>
���mTj�}/�>K� ��
�>ؚB���d�Fn��V�[>�����O���>e1�<=�J�r3o>2�f�%?����+��i��J^¾��>[�q�����|=�N��擼>�?<������L=>���2��=�=���۽f07>?�־F̻�Y�>3�?���7A��@?��޽� K��$��o��H)�=u��� �	<�V=�6��Y�>W%����x����־%L�>�p|������Ts>r�>�b=�f5?���>�+-�&����9ž4����Vq=>��>k�����c�Kt=/l�>I�>��X=�(	�0S�?�|=���i���iT?�G�=[��B >�d�>��>/�����->
��̈?�L���=Ґ�>^k=%Xӽ�	��'oнR���#����N?'���g?���"?�ӹ>�]����=r�7�?�4�=�����U>C6T?i+��d�Ƚ-���E��>?��>�fýL� >?)L�Z?pH�GR�')?N,��:�2���"�@:B?��K��t��1΂>�K�>K/�=��C�!)�=�#��s�r?�O ���>UF�>W�h���>�[�=�'JE>�M?>:Q!�t���B�=��1>������`;�2#���?�2�;�9��1L>�z�=�n��$>�K+��:�>Q�>�zL>ǲ��o/�>Ƥg>Q��=��Ӿ�����>�,ؾ.��V"�]-w��*<����~���g=޲�������h��>Շ��j���9�e��>��9?wJ`=2�?O�V>e''= }"?jS'�Ԟv��j�tű>�&���,�=�)��}H�>�@�<?���{����?�>���E��to��'�9e�>�&{��L���[���j��j�=��ܾ����T�ĢA?g��>�,N�Ng���2w��������Z[I=g�Z=��&�_w����;/�?��-���=ؼ辅؆�|Q?�l��5�L�ܥ�>派�٨>��?==���l��>��r����������8$?� �>�ڴ>��r��<�����>c�n>ڼ=;@�&�d��>�}E�UU�=V��$
?c���0=��ܽ��>��9?Y�'��
>C ؾ㖣��w�>��F����B�>��/�9� >D0���V��D��5p�����;=\�8�Z�y>q�A>G�>�2?Bڄ��!���QS>���>��<݃�<p	�u�!�-�>�uJ�Ǿ=A^�=�o(>ܒ�>/o��]>�b��[� ��H�O�=�n�>�*���]>�����>�F�[�C�J��;Q?8>PJ�=j��>շ�>V�b�^��c��>:��>\�E;�{����?󿾎������W)̽T>�FY<�C�>Ӏ��]��<-Q?!�P=�� >8Z�>tM�>�H>a`g�����RľD
����1׾n�s>�}5?��I>ğ0���=>5�>�3�>�E����>�R=qPc?0����(��'�>�U�>#/��5�>Y��>_��k �w6H>�R��s}>V\�;t=�C�R����>?�7�x`�>��̾�z �h��=���>]�>ￄ>���Ϛ=�>н!�T����>� �I�;�町>��>�-&�HP�=��&�W>&/�>��U�X����&=�Ϝ�֔���)����>@_��?��=�?�z?7a�>s��>+r]>��>\n���	?V"���R=�\?�A̾��ٽ���>�4 ?{�k�Pbu?v�t�\ޝ>������}��<1��>7� ��Q>�ɽZ�?j��f��>�/=�Ag��O>�� �������ɾJ���#m��>x=�f4�o7>����g>��>ԓ�>�%����"#&>U˶>�u���X�=�Ⱦh�>+���?g���>��V=,5�>���=H��>T'?F2�E�=�j�=p�>�6�7o�>�k��'a�=�6�M�<�)?*�^��oF���>���>���<d>��_Y�=�$�t�z?�����>*��>H$�=�L">�Kݾ÷�=f�:�-��w��/>=�>�c�DR=??�#���">�Mཆ����$=�Ե����=;[����.�=���>��?�5'U��컅3>���v�=�����8?�C��������k�.8g��6o=QE3�G�4��E>s�׾��>������>>J��'��DW�W�A=�?�M� \>-��a/�>����> =�
q�.[��_N��?�F�>e>�轐�>��o>�]'��C��1��=��x��p����j� J�=�CL>`8?�i��L*�>B�3?US>��;1�ͽ�\ �o[W?�w>D�����A���=+׫>�a�������|W��>�2ʽu�w=đ��t?�G��о[�����$>��>��ξ+�e=��y=����i���Y��A�=?cm�i�(>�ћ���J?P'��m|A��W��cD��t=@䞾���>;���]�>Xh�>�*?{��zTR�_-?�,:��=N�/�>��E����>�Z�>phX>M5��9��=�;�>lqM����W�+_>�?�����k;v��j? ]Ἤ˗>ӕ$��vY>�	?�?�=J�h?"�>��=��A>��=��>�\�>�t�>�^	�nn�>��_=u� �g\�=�?>�/>�x��~>>W`>k��=$�>�/W=vH?3B.=v�>q�i�j��yT�����=���<��������e����>V���PܾuY� ?�>'����T锿�1ƽ�b5��7�0S���7��R-����LǾ���=}�>���=���A�h��>|��˖�Ȩ��H$��Hr?Wʁ��y;>��>�G:�j)?C:���v>�2�>��>s��F����e?�%.���<���� I�����G�=�x5=�e��W�<nr�<v�~<.]��DL���A=���غ��m�ƽ�ǻ*�Ͻ�p���@���D��uU<b���4�F_=�	�=�!�=��2�6=ϭI='V�<u��=A�=��;x��<|�5�L!Ҽ&ul<7��<��N=��<�YU=@lP�U->=�U񼡹r=Y��=4J =���R�k�Iz�����ਾ=��<��<�:S=��<�SJ��c�����7����Ǽ���/���K<������;x�y���	��J1=Nw=O�=L�:��<%���찄=4�Z;�O`9�bM<�\�=棽*MD�$=!�V��;�=>c�=f��=T�P=]�f=��W<�E�<]*�=%}������p�<aVp<�5�����r:=����iE@���<�]�������J[���;'��<j�[<'�,�j��=�چ=��`<ov�}��$޽�r��n*Լ�S���	��Ƽ��ײ���� <Et漹L��h"=������Y�
`g���==�9�<h�R<p�ˮ�<2���������w��>Q� �p�&K�¶^=/����G��>zY=�<�i�<9�[<��3���<wud=6w�;��(=;�<|�;<E�<4�[�0^B=�_�=&H<�W���d#�{M����=�Ȁ�� ���鼳,�Єؼ�����q���u��|\=�s���Ľ�ח����=���~����$��Z���R��<͹!=�=[=�o=���;��;��n=���<�=���<mg���	�R궽>��
�I��U=�`=���ۜA=R�;��Ƽל���c;.+�=6��W< ����=�i�=��q�5.j=��<�Y.=���=>��=�̽=*�`=+��<�̕<�(r=(p�<pqK�G�ż�n�$�=2���qԿ<����a�3=��B=On���5M=|h}��u�f��'~Y<�����������i=�~�=  *=�]�=w>�ּ�����U�<��S�i���'P�ƈi���1�}�%�P�½���򫫼�+�W�g<:�Ž���<���=�>�<�<=� �<�N+=�?=%��=����?��;vy�=Pm=���פ�<p���C@=pEJ���/:R_����=�<������<�j�<u�ؼߍ�;�8�='�<��L���q�c.��%_='��<�c�b ���	�0!�Rf�
)�=���О'�� ����<������U�s=��UZ
�ˑͼ�-��IK<���<H�߼jyʻ�
B����=K�P=ڢ��鵽`>�<B�8=���� =
�=vѼ�[8<�s"��	��荻�V��<J#=�4���!;�;(�N=2�=����<�i%=TҎ<Ң��A,�]�Ne3<�A��Ѝ�<s�;��<ʍ@�<�/�=� �=�ä�y`���(=�(���z��/
��A�]����\�<FfJ=�ǹ�*�1�u�M����<�K��ǥ��k�ҼL��=��=�b�=��=��i�;o��нn��^���<�׼���m^���
=��?��.U<E1-=��(=h<��<2J�<���=X�_=��<�Þ��3==��<6�=�7J��0z=�P=@S�=��������[�`P=����C�Ľs8�� ���]:=!��<(٨=Ň�;oW�<�����8=z�3=O�=��t=0HV<��J=Z��;��=�=�||=�*�6<�T�<��\=f�<�)���Ҽy���V�����9�y���<!ᓽ��=c��<jw9�JZc���p��<��!=ɽ��=�|U<�0��E������ c<�=NE"=�>�n��<��;=�^d<!�G<@��xp���?�=X���QU.��!��k��=�*=�fn��u��,�<�Mü"��=a���k�-=+�l=�8=)���<��=�[�=�X�=� �6$�w�+����뽤c�����[V�!������<nw=8x=k@��ZI=j�}<��[�Nk2�6H6��2�=�=�h=�}=24;=\2~<ʕ�<�,g�����*�`��=�#��`�Ž���;2X�9|�<WQ�<F�:��:w�̽�:��Ž*d�����h�:�qg���m�e�<���YvR<E��������=���<��1�����n�&��B��
��?��B6缐ޓ=,p����6=�|<�:J<����;[܃<)@���X�<��=�~�=6��=n�=؋���M����_�< G���|���_�'�R�
I��M��Ҽ�K=�F=ZY0�b��B+��jW��G�<�"X��V5��SK=�лi��|^��.a=`0
�a��=Am]�>XɻsR:�� �<XF<ʪ�"�I��l<z�`�J؈����<����ɯ"��Ӫ��Ţ�+[�Q�<�I�=�w�=|��=���=;'�8fB��������<q��<�n�*����o=��L=.���I|6��l�=�z�=O��=�s���>=~)v=�n�T���E��<*�<+v<����M�N=\��<z���,��ܙ���D[��^�:�`=j��=���м����	<����n�U;O^�<�R�<z򥽓T[�C>�����.=�b�����=�<���`<��5=C�=��fJG=KFt=���=�K��
����+P�Zl�[��Z-�YYJ=��=��6=6�Z��<(�@=��=(����<�-<m�=Rxн��˼��\=��=�Ɲ=]�2<Mr�=�R=��
�BJX�m���ͱ��
��sh�<&�%���?���kƼ�� =~`�<_�<bʂ<�?���=C7�;�/�k����<{q�<X���;���	��;�.�<ٍ���<�>�$,�.�<F�h���׻jN=�n���r�/�T�p'�<V7����7��7�:���=~����=۹N=���=�=;#=�Nu=��<̢����g=�=V=��	�~=�/����
�%:=ȿ=6p=�Y�;�h�!!�;ކ�<R%�>�]= ��M~T<�����=�=9�-��-��+:���$�yۮ��c���r�=�g=jH�=�3�<^F<�6;&�=8��
ܼ>�O<�܀=��x�I��hv;��"(=�M';;��`%g�qg<�j=#��=�Y�;-o�<��<���=Xg�=�b�<�ھ�M>��ˮԼId��V���1u�l�5:���;��#��c��\�<#x����#=z�&=��U<V3��e�+�(�u=�� =��ü�	;ܙJ�؊���-��BD�oMB=M�����?�J�;��Z$=U�j��q��R=�J�;�d��Ye=���=�A�RD:̜=d��=>�2��Qf<�k=�w�%�����=�>�v�Lu��-ߺ�#r��s���|��&ț��V��"e�<�u.<h 2���̼��q�ߨ��ૼ.mf���3=� ��u��&d��!8��D���ss��`��������ڻ����"=·=�\�=v���\�<\��<S��<�;�����<|�=�ڻk����3J=�=}�=����S=ڇ+=`��=�������R�,����1�=FA�<<���<��3=S�>=s:&�,������=~S�.����(��=���<`墽�]���=k}�<(<4F=R�:=�?�<핊;ixG�8=x�QR���"�߷�=�t���k<t_N���D�
��<dń;d)�=�&|��С�R�D�ż=���;Ї׼)�4��D=���=��?=f�x=��=D��=�^�<dIr�@�9���7=��+�������2T=������zS�[>��+=�y���<���=q�=�*�=�W�=�­=���<�&%���}=gK=�b�<T�Z8)�-=�?�<2�g�&Q���c���C��_ٜ:�Է;����3�=�E�<����sἛq�=���=��;c(=ŅR�*.N<z�j��fY������/5��隽;D�����e�w;\�ȼ��;(�<#�����ޢ=�T��<j`;��O��]�����ƽy�̽E�T�<dʽ1d�<ca�<��<B���c�<Y�<(M=^8����=l�R=3B+��s��p�=osM=�0k=C�=��<�ڼܭi�C�&=F�C�Yu�<bz�;��!=�{������ꊺ�Q��1h�>t�>�UM=3��	zU>�{�=��i��>�V(�x�Ͼ�K�����5�>�]>̮�*,���=]�?���>=�=������佊�!=��U>�M�>��> B<��S>�&]�V��>�D�=�^>���>�h�>�&?��ξ'�D�l>�ʢ>��>r�t��}��8�>�l������aa.�ΘQ�3B� �:>�
?V��>�Z�>�/�=aެ���\���b>�~���۾����~�����p0�>�_��aK�>�T=k�>1�.?���=Ҽl�;r�:>�[s?��	�0� ����><fP��a���-Ā>���=�`�>zos>$��>6�˽3�Q>���=Rt�>�P�"�����$���>�
�����>򹹾OL>}�5=�m>
G�>9�%�:k<;�cQ<��>���>t�D��e>3]>��5�Q�s<� 	�K��Kj;�W;�=�۾��*�U!����D>$d�d��+��M��>�f��aؾ�����>�!�>���#�v>x0�>�������GF�2C?:�P>���۴ľ��?��<踾}�����=FJ�>]U��A�A>W(�=2u=�?)�>w
�=�^Ƚci�d���z>�t����~?s웽����Y��*ϯ��B=�܆�;E��	�_�!<��=��Y=��lOP���z��>�,��^��S>��?��r���> �=���>�`>ց������r�=C�l>�?���p��=��Լ8!������t|� f�=E�n�2�4>W�t>fDs> �>
ѧ<͝���t��7{�=l&�W�u�����=�43>��>������>O�<U��>,��>��>!�G�+&#��b@����>8Ы:��K���;��>��J��?�>���E~��r6r>2�Q���>}� ?%i��h0�N߹��{ռ�ְ<y��a��B*�>d� >a��>��v8�>"�>{��>�Ө���'�'5�>��x���@?��>A�=|��=�晿����\>�y��ow$>^�d=khd��=��t>���=t�X�݀�3�#?i9�>�L̾P�����>l��>8VR��m��8��>�6_>uf����>�a�=m��>��z��6����=�+?�#�G�<�$����u��>�����y>
�l>yE �&`V<T����'ξ�l-?״>&I|>�+d�C��>�t�����>������<�)�ý�`��U1���-��r�>楫=)ﾻ��w��}Xa�@�о��3����2�=?��̽#b>�O>Z��>����T������uҾ�V=ȷ>�F���@$���]=)Hp>�?��%������k���?�������{��=A~b�ג����=�n|���?1�k>�>>L�C>���>k�ͽs<��a��A��=Ag���U>��3=�:ǽX�?�ũ=6�r��z� +��q��e��һ1��>�u=l[�>>0�>M㋾B���$�������^]�w�=@�=�w����=��I?�8f>h�<8�C��9>ֈ
���?2��Ob >Y��>�о=�k;2a��?!+>��)����=i&�>�@�>�U���0_>��=q�Y���!��=�Y��>$i�>�����\��E�n>�7�?K�>[��=3Q�=��l��=*>���>Aڃ?D��>�׉<�d<
-�	�l>=�?������D���ž
��>Qƽ8$�=M�g>[XX�K�ѽ�.��lC�ˑ%�8TY=�y?09�=��#�{�>1�>����:Ŋ�Bľ h>�ϗ���}>%��<��>���>��&>	�h�z�:��4���f���B�
���T�<��>���>�Z�u��>&�>z)>c������f6?��=n�?����c�>U�#>M��>�b�a�*��^ʾRҎ�.�����߂%�꺓��0Ǿj�>e��v*�<�6�EL�>�?��>�C� ?�=�ƾLV�>\r��^�����Kb�>煫=3?>�74��q|��x�E9�^�ֽ��>OF�?�j��o���殼Q��=I�/�t��#�{�YĐ��X>�Ă�Z8V��d&��`?���>.��7�I�f�?��R�_��>�t�>%�l@e��½�"�����<b�����۾��>�'?!ˤ>@6u��*a>:r��x%I>V��h�4=���3���e;�m槾c�?^h�>�:�=+�o�����bͨ���r���<�p?2;���r�=�_>A�;�=��_���٪>�m��'��X����?b��=��)��ͥ� �;\m�>c�M�슨�)�x��w?�����m��t5����D?""�>�����>�������B�o>dK��.��L�V<��m>D{�>�J�>��?׋�|�<v�پ���>�?�� z�0��=ׄ?�Tk��&=��9��G>>�@>U�>g :>�74>rU�=�E���ﾾw_�=P����{�M����+��,>��>\h\�g��>sq>2��>�">?��ؾ���Ҡ=+�>��j>�����>���睽��оeI��޾�?�|W>�Sh>/כ�Y�?�tg�e�=  ����=���=���>s�.�Ut�<�b�򣎾������d=%e0>���=�¾��мf4?�̌>,�|�mQ����>���>P�M����t�>,f�=�0>�s?Ѭ��S�X����<A�����:?��?7���S|�>(<�覚��9>�Ѵ�,��=� �>,�&>�&�=��=m�?�?�0O�#�hx>蓾���;4����Y�>�O==cw>� =Uϳ>Ɩu=�=�]��[>����ս_�ؽ�D��񭽗��=��*��/�>VnQ>���>��>��<�a2;��ƾ��[��?� {�Q�!?U�^��Y�>7)B>��_�b�
?W�,?^F���7?����^3>C��>	i�>.��=U���=N\=���=D�Z>���^����dl����>�`x���c��i��]�վ<HV>�i�>�?"_�=L�(���=V�?Z�N?�긾����Rj��?2�d��$��}���=�o�>��>@E�>.�߾���=I�>M��>�&�=9�=���7=�mپۦɽ3��Y޽B����Y�����|@K�C�'��/B����=p�a?���<[h(=�0�=J��>��;i�m��!z�|>��l�.�վ��1���m����S��K�=ݲO>�^�Q�>yO=�>�'u�m�
=FDؾ���=��Mip>9��>���>AI>�O;>����G�F�%0=��i	���J��s��3���>B�]>b ��P��=*��r���h7��!oa�ga����f��\�?���I�>PV?C�6=�E�U�>���p��>�ɼ�[X�s7��������'>*
=u�=4����G�>�Y>�M�>�9f��l�=ព�w�]>�䬾���I@'>)$�>��!=$]߾�v3��?Ca,>�fW�L��<3=�>�B?�U��t���=/b��G>��->gc�>��">%� >���cE~�/+���2w��u0�쑴�١��̹b>�L�>����`��>���>�n�>��U>���Q	G>�t =�I)���|=d4�R�����E�z�O):>�a>�נ��	=a� ���½�	'�$��>���=Pĳ>pK�>'���E�\�=I?��0�pL=���>���>T�>W�>�Im]���E>�:�>E;�=p�e��8��>+��d�ƾ�e����>���>\~����>K<?���>-�??(E@?�+�>�z�>�@q����<K�>w�.��΢>!�>�6��#?m�Ҿ�VH�F7�>�T�>H)�>��=�\�>{,4�W)��Ig�yt�>Xe�=�ۦ>�]u�d܍=~¼��2�q鳾Uˉ>�`�>��>�q��o�\>Pg	��� �O�_��56=r]�=M3ƾ#���V�>0�[>�ؾ�x��꽾wMl��ȼ�G�=�>�~s��޾w��� s)>([?��6���_��->{	�=���>�>�y�>	�?мl�=Y����lQ>_�=k�^>����ڗ;����Ꚁ?�O�Ӿ�eK��Q��xɣ=���s6���(��=�;c�]K�F�=��l=^��;�&��vۤ<H�νm��b炙�?��� �<�Є=$��=fO�̉<�k�<��<��I<�?=.U�=S��<a�2=��=�-��}ȼ3�;6��=�b=G���F*<��=��*�:�69=S��;bۙ�����?ƽ�������.ᬽ��>��=܈�;��;�1*K� �g�� $��f�=���;��;]�A��ar�k�>S<L�v�Ǐ=�vk=��������1H<��>�,�p��i�=y�=2���o-�:@wR;*\ >(M�<]��;r⵹�e> ��=��=�>�=q�=��V���<λ<:�=ʁ(�//�����(d^=�sv=ץ�<�,T;ţ�=�:=�^�<yu=s�]�>k<�=�=��k=��4�6��8 Ǻ�:�<&`s;��ɽ-3S<��ü�x��}�:=zx���n��﻽L!]=N���j5�%vҼ'W>��!��a�9�����1�=
OM�#��<x�ϻ�Ȳ=;j��_�;}�`��=�w��K}�˃;�L��=�T=������v�&> o?<o�!���=��w��
D��,���c$=�$=�M������4$x<�GP=t��כ:���m��&X�����64���=}�;�H�?����>3=�%Խ"d^�����>9P�J%�΢����<wGZ�-�}�.�l�BP1����<��S<��P�l��;ԙ=~v�<�\2��z���x�=▻=��P=�ͽ`M�v�&�eV�=�P=ˬ<�_Q=5}����t�St����a=W��;��b�\�o�
ڼ!=���K�q��=aϕ<v7f=���=M�=5����G=��/<�t,�&��=pw߽{M��愽���&	�<�4��,h=j��=2،����;D��<����Qk�-J�=̟!=Z~];2Iٽٹ<�i�=a��=G���ݜ>���=��<I�нH�]�u�.=��E=��A�A����T��Ԕ�9]�<@p罢F"��o<|��;reʽ��Ӽ���;�E�=t�`����;0D�;rad=�4��2�<���=��>�l=�z�;��k=>Ԋ��M@��v���,[��q�<��F��B��4��=�Η���<�3����=;w��^�Z=雸<9��={�i� qt=�[M=�jY�&�=)ɒ=�y<���(J~=��=��.�\����➽�"-�Zt��g�ܽ96p��ʄ���c�i*C=�(��8t��ڬC<>�F	���*��Ri=��=�j�=~�N=	��=8~�=��Ѽ��<��<� ��Ř�<;J����m��<��<Ά}=��<�S�;ۍ��ׅ=�8=�;�6jؼh:�~�G�GZ8�._:���=Ň�<Rc\�l޽
��?����<�1ɽh�6�����#=u^�Ш�<��=��L�:�4��/=�1�s<*���8#=���=�A�=��=P�>���Of*�������ǽ�����?�y;HS=Im��S
=R�h=��$���N=C�=*�<����팴�.��<�9�;�\�<K�4��˗=k�<��=	]��o31=���=���=�Ͻ�PT<�k�<�R��qA���S/,=��(=�}��*=lt�=���;�ʋ��3�=��#<��\=��G<���=���=v��w�<\��=G=�O�=�s~=��O�t�~=+�	=�`L�$�.=(�(=�~>D�`�|'�n���9�<�Չ��<j!�<Jټ&�^�Z��=��<MJ'=���|�=z�+=e��=!�#�+���E�ޝ��O�=J��<�r�$U��[��;��`�q���!�'W�:G�u�h�?�{����= 9Q�<�m���=Ha=-�x=*w*<H��UR=o�O=���(���$<XZ=����������r�)�B��҉��բ���̽X;W�/ƽ�rc�ǗP=�?�oc������✺���=@Jc�C�\�&�=1c�=Z�j�m�;�ڴ���_�	M�=- ��uP��r/�k�3=D>󽖧���
1���b=d0
;>h'�XK	=��=*�;�yZ<)�d��;j�'0�X<߼��4��~<�S=�t	=^[���`H<\�I=󏁽~}o=L�q<�o��R�~B��5%���c?;��˼�����뇽HM-<��<k������MhE�m�<:��<�n-�Đ�<{�I���/=�1�i�=�0=�]���Z�Ҿ=��+�Acڼ���v����ꚽӃ�$��:N��=,C�:�:��	��5�=�x�Kq<�������=I�T�W��dK��C�=�DM���2��#P<ߏ�<�Yܻ�ν�2���=9�=5�<�慽��$=1<A�J�P���Mݽ�#��3��I�<_�=���=o�>����������D��#�={ޟ�='_�<^��Ʈ=o�=���=��<d)�=��-=�����hK�:�Y��xҼ��x�IOT;���<
&�=��ռ/�h�{p���B�=��4��"X����=/j�=e��=�h�=��>��̽G�=+�J<��=n˦�V�`�V�}�$�=�⯽�۽w�U=�4�<{��=nq�<C�<�Eg��u�=��<��&=��N��&�=�==k;��J��L�缦�b��i��4������w:Լzb<.�~=s�:�<��1����=�2���V<��=�@�=�>�;�W<b=�>2=�=R���1\��u_�:_����j<�`=~Zq�niW����=K��<^3=�ǽ��ż�<n<G7$=69��;��h:����=�'�����;�'���,=&�~�}��:c$��K2=��=G�f<������=���<��x���3���=��}���|��
����!<�8o=ks�~jO9�pE��/,>���<ܫ�<y�q=Ȋ޺�P�F�#=Ζ=�0_=N�!��������E=��ļ��	=�#�U�~;A/C��4���n��K>s�<������V��=�g�~E�_Z��d�Z����:@<�5����C���˼������a���R=�T�<��R=5��=�����<�)=߲=�}��2����^=!�=��L�����,��A=7��=�V=�.R������q=���<���<�M���'=Hը=�b�[g��P%�~ȡ��?��s����d��h<�X �88���=��P=5Њ<��S��2l=D:�=0xB=�vн	5�<@B=8�0��/~��*j���8<Vl��=x�<�=��=�y)=�/�<9�=Q��=���<���=��V:1�l�z��=��=�Z<pÚ<��=\�c�K����u���=%ײ������S���r=�*׼�a��� W<�͹��3��<���Y��<����ۼƫ�gx�;Q���� =�)�;�5��%<���=
w�CxZ��[0�(#�;)��g'�<��=﫣=F��-�P=g7�=�A�=�`�<e����s=�M�;����w����@�a�=�X=sʻ���{=��=�6�=�L�ܓY=h��=%=p=�v������W�M@���=U������;a3�<���;yHͽ{�7��ˋ�e��<����*��n2�-�	=�l�<s�:�ş|='��=��;�x=<<?'�=�q$�l
��Ϫ�z-=;��z���ׂn�+�C=�n@��轼��U�I�u��<�.�<�TH= oM�;���\`O=�d�=0�Լ*狼��=��=��;�,=�ln=�w�=6�-=a�<�a��N��NhI=&9������@Y��S�=;ݷ�iDv���|�
�=ޗ���>4<m�=�>��X=�+�=�gW=ܝ7=��<U؊�O��<���=���JZ�TмZ��=�W�=sC =��=ef>A�t=��=\3�hw>,��;y��u\ƽ'!�=9,(��î��
�7�=�%@� $��Z<�-�=��=��2<Q��)L=6S��>e仄�Y�^>��h���Dg��jL��m������ ��
�����<����v���|��܉�у�<�!J��dx��+�<�N��x~�<�5�={�$=#U�=^��)��..�/�>=R8�=�uU�>6=��'=r��=⺽�A�<C��=�So=E�ὁ��<,9��<k�g>�?m�=>,�=�e�=�rǽ{p%� RZ���E?~�M<��=�V�_����7��'���4f�!�9<��>q�̽У�>�����,�>sݒ��>�w�bb/?"��>�vd?�ޫ>���w��=�nv>�eK����'?���=�r �v�¾�)>��"��J>�)?��	?_F�>���2���վ\"�*��<�h�>���=�zC?7��d��=�$�V��=��?��]J���>�*�>��g����@�]���˲>88>P:?%W7=�����'����>�!>��=��&=r�T? I@��	�|�xWG�M�F��?\��>ڎj?H����Y>������>���>(y�CU���?2�>$Y�<�訽����Z������>����-^��]����!= 
����">��>;w.?�D>�����,���K�0�t=M�߾k�9�زz�	��=��!>�_?�25�����>���-���A���S>C��>��>��ݾZ� ?R壼EC�X�ȼM��>�R:>�EJ�S�W�'7�>�W����^��u ����>���>�$�>-�9��U4=hѶ�ꥼ=U�f�R�=�����/G>�駾iwͼ�_��p�,>�w3�L�Q����� �q���q�=�����Sɾ�ㆽ7>:�1=��~��"���S�=R�]�����S��M�>	�;6���V�r۾^8�>)>��m>������^X>���=|R>�WU?H,? ��;�|��u��қ�l��]�k=&߁>0�=�?X�"��/����X�dF>"Y�=�m}��1���|�>G�8>xL���#��D�����ه�>�t�>(Vv?�)*>�����]�_�>��=,p-�����ƽ�._�>ñ>C�J>R���s�>B�G��Ԁ��uC>�M�=�U`>�tt�r^�=�T=��1���F�e��=��>�T>��s>F�B>;��&!�"1�>M
F��߹�Y���7&ľ�[Ҿ�c�=��>��=�!$���(L�(Z��˽�ݜ����>"E�?:��<G��b_�o�H>�&=>��G���?�_�> 8?6�о���ʺ���c=Ԡ��� ��fb>#n���߁>�6�³K=�ͼ�
����>��m>������پؐ��~ʱ�0q;>�J:#&ڽ��>/���+�~>������>~�� r3��|�>�dl>�{��Z�<���=L�<�5i���x@�{�=����`U�>����>s׵�AS?�g���ھ5,��K�>ߝ[>�J>�d>>0�>� �\���=�y���=�6X>���>5(���.=�oQ>�7�>K2��UC�J9�=���=r][����ZXb�>Ci>�6�DAϽG�����>:=��z��,??`�?>z�����?Fs�L�g��^���A�>�">��3��ȑ=���=�>*z��!+j=(��Ҭ�H��J>���>Δ�>.�}>���>�lq�y�6�x'�����0ᾁ}�=?4�=��>34�֜.?�J�=�>�">�0��q�=$>D�뽟�>���>|6�=P慾f��f�Y?��>�r2���I>E����r&>ؾe��<�`2>�?%��>�V�9�����5?/�>���=~�=<�Y��R?|O�>��>�I�XW!<��@�v�)?ˈ��^
?�c�>T��>t�u=h�|1��+k�@|�>�3�>@o�<�,�>O*��Q/�ǸJ�s��Ba�P�G�sbs>Tu�f?��_�=��C?[��=*�g��!�>��������(|���h>-�>�8�>sh>6�w>2��!)>h1Q=SJܼ:�Y�׬ڼ���=u؈�S-���d>�2>�E���,������>	�z��]�>e����`>�MT=�,Z>V;H�5!?!�?H�?�Q���뉾���cp�?Q�x������d���|��&�=�|�=�&?�"��H��;��=,�p>S��a�˽��>���>NF�>V@�>�)�>�����>#a\���{=������>Z��'�������>��\>�v!��iE<�t?�d��K�4�?TZ��M>�S��>�4����_=��B�lR>
��>�~�>�x��
�{��y�=Ĵ���&�>�=�vҾ������{�_>�>�N����>�[���������=lIU>��
�g�|�ac=ؒ�=�u^>�N;�z2����k>��[>�r���G�2�/=W�>W��<����yp���L>�oq>�d�>c
�b~=�о�T;�
�����>�>"���-v��J�(?���'r=��1��x>�>��?����/ʾ<}��'Qa>�)�9�
���i�E`��`���=��?-#���]�4J���i��ߊm�������y>�?�D>IP=?~�|�EB�=��M��G%?*Ҿ�񼾤Tc�8�>��\>d�D��1>�`�>JC�=y��>�v6>?�(�9'��%��dB>m�->�Yy�ͧ�u��>W[~>A��nċ����� 6־�s�>�]y?9��>[,��;��H��>���=i�v��}��>�>��><�[�������Y���K(?��='�?b؃��?F��=��=�~&�*��=*ڴ>6��>�\>*���J���������������=���>�9�=�j��"����?�-�>Vj��V,>]J�"O�>�/��9m���>�p?A���/4�=S�n>�,���ľ*����K�����-[>���>���=R��<���
d����X�N3==+�)��(��>�K缇��=pQ���YE?�`��롞�	?<�e��>	�!>�z1���&>[�>��ս�>�q��>���=� �=h?�%٥>�>�>X�.�a���ľ]�>خ�>��K?a[�>J8�>�X��tbw���?���B`�>JLY>̵�>����Ύ��X��i�=Y�>>?]?�ؾ�R�=ܼE>ݩ>�`Ž�?�=fc򾩮>�v��
?>�2�=��X�4��F!�\�)��TG����>D�>���>��ƾyQR��fc=���>`0>��=��=�+?�i�4�T�����>����ޗ�O?sS��!u�[�(����=:c罹{�>��>�Z?4n�>Y�x��Z����žhX�R�C��E�����>��
��ؑ�)�= ^I?Ys"��|d��Q>�@��q��d�U����>rg�>��>�e����Wk&>|���!�>QqH�L�'?(rb��s�u��>Q��>�۾;=-�������0H���k�=��>��۽��>U�>,Eu�S���Y��X$�>�f�����=��=R�>z���r���
�Џ8>>H�PC���j�$�$>�z����>!�u��7��:��=���=?J�_�����O�5���LX�>/G����j����<�go�� 9>�Ә=��&?�4����彄V8>ٱ=���ہ>��>�N>�7>/^��>#T����>C1<���g�($�>O#�>�O���j>��?�w�>g�	��풾����Gh�>H�>MK>c���? �=,T�=Z�t�Y�e��f����=���)3>x�=p�w>�x��Fپ��f���C���>;LH����=S]�t_Ž=h⾆�̼SO
?�F߽g��>���=$&�>瓾�|;e�I�q�½�U;=�y�iq�=�iվ�y�;�{���4?$
��[�Ф��f�>�.�=<ٷ�&w_>}C�>M_�>��=�q����=��>m�z<( �+�'��P>(6�����^�ڼN��>j;J����^����L�>�b�=4I�>\�@?�r�=l��>�;>�m
>�K�>��3�Aiƽ�K>�^>�	�>�-[>]�S�0��>5��<J���|5>C8?wm�>N\��A8���\?KD��<�>�y��"_2>iĎ=Ւ����2�O=W��;��l�I{���H>������8�����ؑ?B$��
�kuv�S
>9�� �e?����F��5;�:���Z
��F�>q�=������ؾJ�
>��-?==>�O��>���<�����5'����=�'?��=-F?�Ҷ����=�Gļr�N?�r��k���Đ����>+bc�p��=������>��R����b�7?Q���~�0?S%׾H@O?$r�V�:'�
��>�f��!������EU�����<���=rY�=8>@��=��?�B>�:���� ?�
�?_�2?՞>��>ϛ�>:��?E?�-B�\Jp��v?d7�>�)>I���&��r�5?�=Ǿ�	��[mY?��!?2�D>w?Z�/��^N��ķ���%>=و�L	�=xj=93=ŝh��>��0��0��"|�-��*���t<tq�Xe�?��?�?�ʧ�)�>�=�?i6"�"L1�'f?>�N�=U̽�w��u.>�R?�d�>�!���#�QB�? 2�?�t�����>ڡ?���>C�-�'Jn>�4�?I97>���~�2f:?EH�>̠l�a��><yF?¾���}N����>�"��`�=_b�?_W,?��'>��>{�=yx�>DC���O~=.���K'�C{�>u�������۾��'?E����{�|Z���u>���<��ٿ%��t�?�Z?��(��zt<��F�2��H���Ѧ����>���=��	�����*�>?>
>����)��$4�j��;CI�����}E�>��?�= �w1�w�E����>8���h�#?�k��K.��%<��y�;�Ֆ�M;>��@>�]���R>�H5=�������[?�i�s�ɾơ�����=�	�Q࿾�-Կ�~>�gB?¼b�I���v�{����3y>��!?x��������>�?N"b>�	�=y\�?�Q�>vI��ꝿY���F���&W=���=�":?�l><��}?�
����=�+?.z��2V���o��㞿A�v��|�?4�>���> �>,7!>��?���>��x=��e���I?��A?j�%���n�Rs�>P���v/��Od ���8?�#j?�.W�Md0?��y?��ʾ7mK?��4�CΠ�G�>�J�>�.����u~1�,��=���?n˽>�W�>7����o��I�^�	?���^c=?�I��u��{�>&�>��
>p��=L���q���9���=�L(��m��� ��b??Y3��Ó�V���ܢ?q��ȕa�Ǆ�>�=�?�J+��v@�9X1�d�>������>?#�>��->G����� ?��J?������H�g���z>��F�h��=N�??l�g�𿊾�m.����
��>�qG?���H0��?Ð�?#@t���1���8��Q�>j���{"����S>���lk�PÖ>���>|?͜��u?�?�Oվo��j�D����>T`4>�8�>�nE?�����Ml�ľj�S���q\0�tͱ�T�?<���Q���t?��?��弴�=��9?�B:�!,>zE����>� ?��"������ٿ%?�GA��i��(����?�ֵ<��x>YN�>E���	�ۤ/��?�s�>����3���?������`�~,��f>��ྔO�[���?}DT?�?�*?h�D>���>n㣾+n���_?��������n�3?#n>gY?�؀�����t:��X<�a>��?�i�>\ɹ�ޑ?���?F��=ENS�����k*@��m�[U��2</E�?�D>;�|��P�>Z��?�y�[�-���[�ي���dK?��>�'g� �`?��-��d�>3=?��c�:{�>Iτ?�9?D�f?�v׾V~>���?�����>*� ?< .?�;��ߍ�=�P����&���aȇ�#�?lWA>:N>!<	>�01?:;Y��A"?H�>�<7V��]�{ī>��H?�ا=U��=m��<+�?��?���>"<�=7j��r1?���*`=O⡾��ﾎT���-��fB���><�?�K?{]N>�ө��
�>p���G·��tv�
/�>q.?u�|��w���?�ʾ?�`!>�9�������=����\��@>�0��2��_�>|�澰��>$c����?�N׾�C����V�+沽y������R�ؾe�?�|�>���>��B�:-���+?���?7_���� 8:? �?΄���0�����>�.�?gD�����~�>�Ȝ�G
��`u>"��Wn�ˆ??i�4?	��Z��6��>)�?t���DM#>ou���?$����xS������=���42����>q�?E�@?u;O>�Y!��W��Uo��/�9?��S�D�W��>�㷼# �� P��s�;>҇ɿm�*?]A�=l�1=��>Y�g�Q���/7�.��?a1�?���+[Ҿ^]%�ձ?��?����5�?:Xm?�̓�(r��뷕?�gU>xT��>O��P>���wN���RO��� ���>����F��n���:#(�����;Ǒ���X�W���њ��ʎH>h����>��n?_ܽ�򾋝u���x=�x���J�9e�>rϣ>�ֱ��C�$��?^��>efW=�1\�nks?"�����?DԾ��=?J�=[�
?�pK�0�>��c����=�#@?��C?5��>}�.���`?�>�D?�e��ھ�:?�}�J8��ʀ��@�?䷥?ۓ��h�?�[��J���*�����=��[��t�>f,?ҥþq*���ڪ>1_
?���>;顾y膿''�o�t9����qb��u��ˊ�=-[�?\=�"���_=�"�?��>ՖҾO`�>�ͪ?���o����>�qK?S�v=&����xC�5�=��E���׾�&���-��Ƞ<��ǩ����%�3Gվ�jʽ���j�>\	>?旾��>KYb?��<�� ���:3>��?�a�V_Ϳ���>�P?�~��	)���ľ�d�>	jn>ټ ��y����=#��>�d<I�?�t�>�wK��閿�h��(�>I^> �G?H2�>D ?��> �>�뒾Y�v?��?0н�(�]=��=��=`H�?�
 ?�"V��ޟ?���M�G>\˗��
>U�+>�y>���>B�?���T�~ ?dȽS����0>4	?�纾vоJ:��6Ql��V;~0-?zѐ= �Z>�SF?"�?j�����>,�"?�{��$@���@��� ?��?�*�ZΌ>?�%?�*=��'?����Ǧ%>�8���=��]>��=�uU�A��>�V��3?�^T>�����_V�r�U�Ω>�r�>�^>�?������U?R��>?��G�3�B��
[>�e�?��>ں>�_>�<?!ô�����4�v��U��>ʱ3�/����X�>��~'��`�j��lD>�?>̵?�E�?[�=�����w��ZL���>˘�bå��Q���8�>���V���
e�L�վz����>�F��<��xX����?.��C.�d�ľ��{��љ?�?��=�ܢ=_�4>�y����g={%���=����D+>~�F��rp�[l>��?�	A�K�۾���M��?v�>�=�>��?��K��<�����ࡿ���>��>{-����ھ�?�U?2�>��$>�i�>-Z?�����L�-�?>�*�?�,��\<ܾś���ٟ�jo�>����3�!�����U=��uE��G�C�.�ƾ�#�0�u�*y4�Q"O��>i�q~辫�n>�q���ݶ=j<>Ӽ���>���ɾ�uE��R#����$~�ͦ¿�`�>�	�����?�	V>�A侞���x~W��Y������0�� �?�f`�<�K��8�>�?'��=>�%?�=?�O���O�<y���@�*^�>b�<8˽%'��J�� s�>�#0?�%F=�@?��s?�6?GL�?͊9?v+,���*?��7>DU>Dt�?�Ղ?ݓ>3�E?r~<���0>Z/[�!|W�ӟ?v�x?4ﾹ,��d�=#�9�Ԑ4�t��>A�?Ok��ݹ����z����>�P���Ͽ�Q>a��Q���K�<���z>��=E���)�����?�Z�;�c����t�R�|��sN��K���ľ�ϾK䪾BZ������V��=4FK?�C�=���ၱ?�!���b���!��p����$?�V�>x�?!_>2��>M��3�?��<[t��Ȅ���	?^W >��(�u�q?ŧ?p�>ȑ������Ь=A�f=I1?�ow�k���v��>��j�F���ݾ�ľ8 �>x��X�d=v���jb�>Gܘ�)=J��e���-�>��i?�|>�,8>�>?����:?��K?�a"?}�?�����!4>�?K!?ƐP>��>2�>�D�<t�ཪy =.(�<!:>�X�>X�>掽�"&�9��V4>>�N��݉��ﾎ9\?�R�>'�m3���2�є��`/&>$2ξHc������A?^���6�m?�)P���t���r?$�>|S�����T6_���'��"-?�j��l�˽�c�>c�>uB�=���>։?@5�=����Y?;��?$�W?HhY��Hh�8>z���?Φ���@�OǦ��M}?��b�N�<y~�bi�>4%,��?�OPW?(0�!��>G�>�6n?Z�4��8=>�h�>9i�O6��� >���>�zQ��׾l塾�����	����(p���#Y��x0��,?\3?�y=M����i��sU�=4~P?�,@���,=>��>��N�:�7ߙ�� \��΂���:�..�>s���AI��a�a�z|>�e?�6c�S�-�!ਾ��7�}#�� ��=K\�j�/������^���=~L�>]���ý���pw��З;�i�>��ξ�f����s ��9��� ������>�>'� o*��ʇ�V!�>�G�<�z��JJ7�P+� ��>mQ��u���\�H�F��G=<_����]��a�>�c�>za�u���iT�dL��db������4'> dA�p��>!3"�"���F����>0�z�3��=�C�){>��n�R��>:C�f�>�a�=�g��v�̾}K�>�=x}3�[R���ʓ>~=��\ZC���ľ��.>�/�>���<B׾Hf��z�>�`�=D{I�c�t?㾼E��� ���6\?��ѾP�ὧL+��j?��>Ǚ?Wd>s�7?1�'?��?�r�?��=^GƿpuQ�|��$c�>k|���׽�� %���H׿�r>f�6�s1?�W�[)P>U�$?!]1>x5�C �=���,t>NB��h^�>攮>�8e�������=�.?ٛ,���">D#�2uO�#oC�a�佻ʾ��J���(=;��;�7>n��<n���*<ľ[����w�>ׁ>]J���>EN�,eo?�H�>�D�?�h|���?���H�?�y��{2�=���V}>������[�O?[�?p�?�fc��6�>� Z��32?�A�=��<?_
���09?�N��2}.�֊�>)�!?or��g��m�??KO�>+��;�W�U�?H<<��Be=�C�=�"��@�.�����7?��B��v�=ƅپy�=�\5���)?�佸>�?C|D�=�>�R�<p?�3׿`�����T�lrܾ�%�+�x>l�?��־��>���9�ܾMƎ�+�?����|'�d���u^?!��>�����fX>J>?��(��6?�b�?��q=91>�b?��>��A6�Z l?�$�?������	� @?q�W?�ؑ�+�
=Y:�>�C�>?��>�Au>�z?�8?�O^>-]�=A��<`�$>��A>ړ�ɛ�>�!�<�g}��Q?��>ة����@?^؅?0�5��?��_�Ʃ3?|�>���:;�>"]?� g?%�a>'z=���?��$@0f?q��>N˓��̃�3�q?��a��̌���> 6��w�>2?�7?��;.=!?:��?}6>Q�D?ݲ�:%�j?\[�>��}?�1)>�^?���=�p?������>���>�U@�Gp]>�P|��|�>+#�0?9�S3�N��D_m��
>`��Ͼg螾1C?V�9���=,7���f�`7��֌���?�QH?D��>������=�Hv���?�!�m��>R�??^ =SL��=><���u����&��Q??���>��s?�g��?�(�>�my?m(� ��>�f�m�u?�s�;`�z�b׍>�������q�<��!�7��̛>�?���ھ|����'>?������=^?b�)�¾��o>��>�ˌ�}
��փr?Ồ���ž�;9=^�?�/�>u^��%K�lu�=�y��S��>�8�>c@{��ґ��9��R`;��08?��q>��]?��"��i�>2�>�*?�L��R�1>�_����5�栿.��0?Z��?�M)?�4�C�������ZY���Ǿ��꿲gA�H�/?�G;��Nu���Z�=	���v��7��>�c�>�����Ѿ�F;�ɨ�>U��t�<��ұ>-��>Ԗr���ξ���=[���aN���><_ҿ=�5�j�>�>!!�(�>�A�>���s�?�ˑ��B`Ѿ�����I>���x;�>(�7?w7�?Ϩ=�r��h��w-i?ؕM�i�(���n��(9?���=��>X�0��G? �a>��?3Xb�D��YKX��[���;z����= ����Z>U�{�E>Fއ��s>����r�`1�?�{v?f?L�?�¼��F���>Q�,>ֿ�蠟�ȇY������!f�=����cRξ]O��9#l?�q�?��I�g��>��>&e��{��6/�����>�[���C�*/�l%<>��ɾ� H��ǝ?ܷ�?��?��G�%3�=�Zs?�#?oVU��t�>'N�>�F���]��2���Iy?ͦ�>�(ý�e�>�@�=,�C������󾯢x��"�=\
��>�+���=���J&�=��J�~d�>�B��F
P��^ʾ�6�?1���ٛ�=�_����?�����ﾮ�:��[? ,<J�>4�X�K?��X>Ȗ!���-��L	�	˾��>F��%Ȝ���%>lF>��>d�w>�?�������>>B?I�=�T<�y?���?j�x?c�),�>M7?�K�j�<�#����Q��?V=���>uy����>��?#��>���nK?�Od�ଛ>�{����1�X���p��+����>D+s���� ����c�[�?_,�?.u>�&^�ۘ��L�C�
?�6Ǿ�P�>�}�>�1;�7�=�ς>��?$�B=P�+<^d!?u1�?�Z�ח��B���&�?����0��q!?)�3��V�>�<��z��>�y�>������>�%�>�M?oy��F�s>��:>��?F��=v,?�;�=n��>I�=��?#b]���>�>��:�v�>#C�?��T�k6H��h�>-IO?I�>B�>�o>/�;?ʋ����6=9>����p?���_ݼq�=�h��\��>x�E���'�	ط��CT�,
���,4=�/�}�
��m�a>?l�+�������>+����U�$�N��>+(�>��?���­=Ъ�>�],<@R�@]��a�>)���z(�m6?�@�;��>$�&�M|�>���>y��?ʹe�X(�?)�a�;��?�ǹ�zz�<�}��,b�>pY���>�?��0?��]��
$��Lʽ��e<$��>9���5�>x�&�'k�>?�1��;>���>�>�}��.=�Ő@�K��=I���c=<5���B-�S!����)�u[�C!n�F����]>>�����<�c�M?;�/��e���ٽ�^�#b��M���lž�>F�䐬���Ծ[(�=��{�>�>�<V���ؾ3D�g=?,�:�\�?��<�n�ž�X���2�	��oϮ>!����}?qz��@��=��>�>Gy��hT>
��!W�>���(�s>%�ۿ��������U��f,��9�L�_žl��>�t`>`���Ǟ>��<K�>�J�? �y?g�>�?>��*���>䍇�����Vz>�R?��)��B�>�*"���><�>A_����>�Ǣ?:���U�B����Q�>*hӾ:'����R�	 �?��L=;��=��=�?`L�5Q���B7��ȿ�����E��n��~5�I6���q��˖�^熾��5>�N�K�6��l�HK�0�y�gb��W��>��x>�l�=���>�+<��u?��>&�������>��^?�B>���%,�>�RD��?Ⱦ�Q_���o��&?:H�����!���Q��UNŽ��0�I�=R�>�a��|�<J�3?���>�	���=w�&=�J�����9�?3�=.d��yw��Y̾�S�6"��2�A�=�¤�,�>��U>�_���_?��?�B^?F݊>G�����>�?��>��>g=>ԓ�>�σ����=��=^�1���>I+<P�>�s�=��z<�Z?p�>W�����G���ݾ^4о�S޾U�T�d��>��>�3�>d��>[]۽����E���?ƺ;�m��Cu��I�������	��*���T�>�.㽵Ŵ�g�#?V$�F��a>@�6?�}��O>��<YS�>3?)�DFC��1~��ƙ>ۛ=���>��?�y{?<�i=(�5>�Q>��?A��>٣�<+0�=I�W>�U�iR���5�=���>��=���1	������tf�=�>yZ>l��<}����4?E
�>^ɽ����JUȾG4=�>ɾ��¼H�=�����s(��ϕs�W������S��>b�;�?���^��-�>^p�f?T�$�q	��A�>����3�&��$$?�G><���eپ��P?4���L�ܽ��8��L�>8�D�j�e>��=C�]����>w��>GT����\?�_����/������Y���>�̫=�y�<z�>�7��D�ܾ��)�j>��|>[4��M�[* ���J�'"��&N�>:-F���*�a����6�>�3+��G�=žU���X��=T^�=��9�����B��8�>t��={��V��>Eq>�a�>?	:������:վ�M���=�̋>��>߽�>n/�=j2�����,���̮>z}N=^��YA�<�և>�ꐾ�w*=�(">�����>�W)?�@?�؍>�S�>�L���2Ҿg�I=�7���^ﾦ��$�=��ܽem��<��=%��>�i�>�-�����>L�?�"�=�ݾ��3�!^�>��^�F�V�Vd��E�E?��!>9�>��>%R5?`@�>����0��޶�������>B!��ӝ>���>�x�==�N�m�����Ծ�!��c��u\�{D����
�7�>!�5��A�=���>��$?�Vl��� >���>C0?��̾�p���->Nz�>���>34强6���\�/����������q?�ؾ`�w���ýa8>�>��������S']��Y����>d��>|�Z��>ܓ�>Z݂>�F��s=�`>���>d��Y��$>��(���� ��8�þit��P�?���M�Ҿ��b��o?���`t�j��[??��^>�A^�bթ>���>]`+�A?���F>�?�Þƽ�N,��	:�N	��۳�5�#=�%�>\�ν�{�к>�c�<��"��r�������=�iվ�'�ikr>��ѽ�j���>@�w��}=κ��ҧ����y�����>�~">Ǟ齨7�>��>��ɽ`Ǿ$�D=�ޛ>��Zʽ�>-tf?)3�>��>���>o���r���侓���4�
�cL�"��>@?I�[��	�=j�>i%>=s�>o�<��>�(>���=-ɕ��U�g�?A��q��=�T�=]��>���e}=�BN>ɷ�>7�[�ȃ�>�%�=�Dp>���~z������������!��v�>\��>%�� ي�/��>
�?H��>���=���=j�>��D?f�>��D��'���yD�tQ��W��>�> ?�=#s�`5�=}|=�B���rT�2������.�i�������N��P�>�=ѾT�#>8�>��>6U���g�>'�D>G�\>'"㾹��>VF(=�=h�>i+�>^.�=k����=�u��Tݽ>
��Z�>�t�Qw��Fջ�S?e*d�m�>��>;�U>�a>z辻!N�YM�>/�>�m�>�+� �r>�/?�ފ>F������9j�gq������q�{���M۾i�L�75�.?�<pw�=Q���|mƾ���"C=�E̽T� >�`�>�l�=W�n������ξ���>1M�?�>���>�yX�>�����#��4?��.�=̦�=DI�>��<���;�I�*RV�d�����=��=BC���3=�>�<�����fU���j>���>M5þ $�=%�ٽ7Ĳ�}�v��g�=:/���s�V�Ӿ�.�꼍��'�=6ҟ��<	>QV�>���xk���cN>¸q=����Ch>�V�>��n>�ܨ�C�ؾ���>�^4>�=c�|���{k�F`�͏T>����##>ԧ�>'� ?�C�ʹ6?�q"�	QϾ ,���n?ِO>�A��������>#��>oG�=�GݾP�>l�>�ꗾc��o�߾�7B�eԓ>�~�I�;�w>�O��1ѽ�-���Z:����~?��'N{=��>A��>�46?u��>��>5�
�v��=kܻ4z
��<���>(�>ry&�Jh=�>�(>�>�!�>�o&>�:�=Diӽ 2�'ځ=C��>e��=�O��]�+��(�=�b辁�����C�w=P�c<֛�>�|C=H[�>�a־J�t��2�=�1�΃��B�<�%�=��ľ�1d��b'�)	վ��>�7�>\wk>w�;���=�5>2Ҟ������6�=�c�>b�=>ޛj��d���پ9��]�:��@I���s�W!���;?1����@x<�J>_?��
�D}K>m�{> r?�E���n�>�3�>��<?�?��ڼe	���������"�o+�>��?r�m>��??�4�3�˾�\��\ֳ���/�8=�.>`lཔ�0�kp?����V>u��C�#�=��=��5�ip���y$>��>��޽�>�?�>���<2�|,�=��R>zZ½e�ʽ��=Z���w@�>#꾕޺�̴^�P�?"7�>r�\>bf�>)�ʾX��>���>*o?���>�$�>D�A>�=N=�V�9�`>+ky=QAM?`>�>�=�b�>%�?>N>������K�^�}?г>������-��.>Fg�>��9>��[�����c��?����s�&Xr>{Z!�v�)��gB?E���ә�= b�>~EC?]_|���9>Ć��)?Y��3��^UνR��>@?�;�!���=�n6��H>X5>%c+>h��=[��=��$?�s> ����p����ȼ�N��!?��0&��~��d��>��˾�N]>��>�G]>�߫���>��J>��>m� �eg? �o>e�9>��A�>&�Q�~>U����rm���U=�|��N�Y>��H�K��>c�=g�u=�k��� �>8$>ʕ��-�=��/?�}z>��t�9��>�:������B�>xq����W��CT��!>�#�"�a뉾��;�Ż��$ƾ�;D�X}G���,���=N�Ƚ�.��Hͼc�<�6���>t��>�Y�Ȓ�0����w�߽�q���)��~>7�>��Z�����GeN�q�>5���>tϽPÝ>?�=�OK����8��7Ѽ�o?��7���=�Л>R�>}�%���=2�>A\X?An�{��>乀�Q��=ȝ9>�O�>��>-��s�>,(k������X�#�>A*���J�gZڽ�r�>qC����W/Ѽ�3�<;�?J0�>�?��� [>�;�W�F�RzI�Mo<?�Й��"���]��8�0�}5g�S1�˵f������Ǿ)�H?Q�#�,D�;��>�#�>�M<����Q�����?�Ȉ��߆�31>Lz�>�Ƚ>4ݖ>��= ���&O?^�$��4]�2��'ߟ>x�o���Q�J�ؾ��?��˽�|=L	>�S�<�8%?��>n�%?��?+ *?cI>��wӾ:��>/k\�U���La=\~�>P�d��_м*XC>#��=/o?ȍ:?S����E?���>t嗾G�^�1~�>i��T�;eؾ����0|U���	���I�P�B=Җ>��>c}	�j��>�+�<�j��E����>h5żE53����Fᙼ��׾�B����6�0��`�=ޟ�!m������$>�.�=~�f�"�̽O�4>���=�߾h:�<+�=
�=�>�����W�W,�>��?c�x�W�q���=��Ὢ
��2~�������>��8tľ%
ɾ^��=YpI=��8;i?-�8Kἆ�j=m�F�����9����B =JB<��%�7�A��I���<├���'�Y~d=��2<�=I!�=��8(2�=TXU=��=�!�6�<8�#<(6=��=�@793�`=�.:=Dk��b=ۂ�=���k~�*�=6�M=b}�=%��;�Z	��$<%b�;�F�:u!點����� <ؼ:O�y��<$�<��c<�Ἕ���@,�<��;%>=�>6=>f��+�<RO�=;й�q�p��hI�Ҝ�� j/=��=�蔽4a=H�=Y��=q���<�`�<:��<�̑:Y&]�������=�8�=�]�=@��=]��=��޽�;;��HJ�=XY����<�-
=s1Q=Do>���;j�=�$$<A_T<	H�=���;M�c�Tv�=u�<�>p�U��럼�B[�6,�<�7��B����̽�����[�+�t���7[c��pϽB��=��M��j�%^=�@9�=H\����=��Ͻ���=������<5��Mz!=q�S�"��MX�i{
=Oy�<���2���J_7=��ҽe. ��'�̒�=n'��m���g�\Ψ;��=F"�s��*�=�f�C3q�JZH��u=bွ�J�cx)�+7��|h<F�>�QT�+w:�E�&�h�4ѐ��z�=+wZ��9X��N�=�x�<�����S���0=Wl=ur�B9�������=L���$��A�;�~=��=h�������'����='G��h���{�2 ����ٍ=Fz{��&=�N��h�i���<�A��#+�[D�Τ��t�ܽ�a߼�^�<�=����=4��Wc=�^�c�<=��=5�����G<��'k:�����2|-���;��<��v=(z>q�@��^��Uo>&9?�X;1=��6=p�<�p3<T�"�8�%�yq��;T>�������=�´;�8�=��=T>��<��=	zN=��h�<�`����N=u��v�<�w�<�F;��.��ڽ�3��8Ɔ��ս����b����=(�<����4>�� >+q�=�sȽi��=#W
>W�=m�>�$w$�j�=>�=Ѝ��c༈��>o�;�f"=�k�&Y��_m<�����<$���=ѝ<~]�9��G=Mʼsi�=v�4<h�=H�$�,����=@��=��#=Bs���)k=�'�<H��=ދ��%�<莽!�o������=7_ü�P<<"�'>��ؽ��^��ͽPN=d9=�:н@�=IQ<LP=�}N=��)>��6>�;��=oX�"�ڽ�T=h�ѻ��W=ƭ���MS��|<i=+�;	�!�]���p�=�!&��~�<Id�<�@��Ώ�<O
��8�=D�>�፼��<p�=8x��w�:���ڽh�G���;��=�竽�5�=��=��!��ƽ���?2=v1�;�Ц��F��tA�=9��<0�=똧=kj�=�
�<�O�<#�o�h�Y��=��(=��O�)ə=������=��<cp�'^�<b!���=ҵ~��u�>�=3��=��=�j
��	6=��=�]>=����1�:= C=�w�=�����Xɽ{��=���=��m��V=Ԫƻ'm�=�H�=�2I�1��=޶ݼ�B����Q<|����xu.=�P=3��`���\�f�r;r�*=���=����$�=��ͼ�x%=��J���L0d<���<�]^=�{ �2����\<��n���4='�4����=Q"����O=R">��=�"��'�=,��=�=����ɒ��߀<A��=�y=F���gI�����e<>��<���@�;�+<�) �h�BJ��.<B�=>Ӳ��<��@���C��.�����=��=8V=��m���=�V>! ���s���#�<4����Bٽ��@��aq��~�����|����r�=�=��;�MK�PJ��H����%мZM���=1t; ����<0s���/<1D=� .�n|��v�M�1E����奕�����m�=&Nb�n��=������w=�B��yI��`߽�����#>��Q��$���>=�ͼ���;ƍ<uS����Ի��<�%�=R�ż�W�;K����K��N���v{=Oc�9��0���(��;�1Z<�ֽ�P����<_W����=����ʐ}���}��M�����	���*>H\�5g���
��Qlʼ�(��Dܽ���q���m#�<mg�F,�=�����ֽ ���(��<��	��=��8-���Y�=S�ϻ�#��|��di7<��=���A���|�)3���� 5ན�����<�<�=�#i�n==1v��Ǽ������ޞ��S���:�:=�H=��>�>B;��Y��n.��(�;,��;���;�g$��p6=зN��=��F=�=6e�=�I��O�O=���)<*<�a��ڛѽ-\�=1]����=��;��F<��"�!����H��[�������=F�=�3=�#�8�ܽf�<�g�<���Z�ؽ(�=9��=8B��Hf�Z�]�=�q�=�i=���W;�`��=��";B��;�c��7���iy=t��;��J�/B�����*V��&~$�L���	o=���=��=%B��
�=�	�=�^�=P��PT�=���=��=)���ʑ����=�i�=��M��!;{�f��Ƚ��ͽ12��cE�lWn=���<���;��l=1an�����KQ�g&L�D���\���H���M=���=�7��_qE�R0��0�<����Mjt�k�ƽ�J�<A�ī�=3O�=���=�SU=	���;��=8��;���j���*��=Ѹ��%Y���X�Z��=GSz�'o>�ω=�=��S=ly�%�q=�=���s��=�ѺG{��X��=�=`����<qBM��@,<���*];����K��:�}�=��<*Q��C="�)��?=k-��L�H�� �g<b4��JR��~뼧���T�=S�=� >�>Z��<�'�<��2=|�=��ż:=�z�=p-�=CO�J2o<훅=ZV�=?@^�1J=}���O��nP�������=A�<e�0=Vs���>��X=$���H��]�p����<���;�&e=z�?�n�=5��=h�/=S��;��<\T�=�a�=�F��b:k=,P�=u=��޽v�=������:��4=����&�D=R�$=�U�<�+ͼT��<�E9F�0�c�?����P���Eŕ=��4U������=�偽�0��Cm�;�$�D���C��&����ǼaN<�k������M=�|`��F�o�[�����ɓ[��/=*�=Q�,7��BFn�9_$=�0�F,༡c���;i�3<�=؊¼E�����=�9��U��=��:��=2�:��:����f玻تr���=O�8�Ѽ�;4����=��!=�3�!'>�)=��`=M��:@r=gT=���=�����������;�FF=m.d=��Ѽ�N��}n�5uӸ9�|��{��a$�#߼O�n{��hƼ�����ľ:�L�*Қ�<^��m������=��=l	��({�g8�<�:3�������V���`<�BY���ʼ��a�k,��M=��W���t�=�g��s���)�_���kV�����툓�q��������<0v�=^r�=p��=V�8;W{н�y��e8�=���n��}+v<m
���&���Ƚ5k���21=��=-!��Z�����=�^Ǽ<�=R:�<�y�=���=I$��' ���)���ak=e]�<�n<�M=uq�=�hY=��;��#>wU�=7||=%��<���=������ͽ'��Y��<A���㡷�h�Ѽ�O=�f;
xC;�������<<Ч��ݴ�\1ֽu��<ߗ��]��3���W�;�?޽%�߽��轈�=�����ͽ�!�{Q3��z��޹P������k�=���=�z�=D<�<_,�=�5�<��k=[üU�=Ԅ�<��� g;�c�b(��s���A=�/ͽ(����.m=դ�=����Q0= 0���D=8۽Ck���A=�m�;c�<?#�w�JzS��'O?���vu�O�~=��a>�̾��j���Y���y��g�9����������>c��>��?�/�?��L>���?%��=�?��= ]�>�ϥ>�W?78�>h��>�9?CZ=?s@.?�#����>.%>�.
?���z��?��D<\`.?��U?�V��Ӻ���/�.���ؾ�m)�Q�><V{y?ǯG���?o����]Ͻ`z>�7H?�\�����>K��<�{�>.C/�&�e���4>�*����?�g*?�s<��p�[���ű�=�9�>�}��{���&w�~dV?\�'�QO0>�?����]�=5@�M�>0��?�A�����=@�#?�O�?\ڂ�Ger�D�>dw�>�z���'�0;[����>�=�P�Z�[�?��{׶=ӿ=s�A?ڽt��H�>��J?A��bS5�k���$ھ݅=��
�4Ě>�>w�g���K�>�?,��D]�� /�Ad)��@!?��C>Skݽ�>QlF?H^0=��?�<<ԡ��kDH��쟾��<�!u��e���>�N.?/?��R��D�n�w?<�>cK}��U��/4��{�����u?(���2�>X�<��L�\�o�j����-=8�e������,���Ⱦ��6>.8�(�k>��*�����1zV=�4f=�d�����0a>�t�֔���xv��K���c?T�"��Ѿ�!����&��	��d$�?����|u���m?�^	>[T�>vĤ��a����> >�=����PI��M���I����A?)D�_��?&�	�XS��H<B�$?�2�<�e񾖞x;!�_4�>Cσ�jW���?T�d>�3�?=O�=J�?����*�ྵ_�>�Q�>·���P#��T׽!��!�=V�E���W�{���<��B�>��C���3?��>o[�^*0���'?3��>E-�$S׼5T"?�OM?�C?H_�=��
?��,?�S�> ����>��0>�\��pV��?B�>���D��ud�:h=�A2�AW���7�>D���Zg�i?q!>�]��
�?i�P>ݴo���t���s>��>8�L?�3���$�>̥:>�舾����n�li;>9ߦ�A����qz>I�� ��޼��G<�Ys�m��_�!�HP���>�
U��Q6?��6�ǋ>/�*��A�>�n>�3�>�`��w���?� ?���>I����F��r��dnq?�����$S�I4?����@?��`�!t���6G>���>��پ]d�>�#�=��J?؃�>Ѯ/?rԾ��A?��>��������U)�p�?����@??Ĉ��:�?�]�G?�?�X)�J�>9��=���RqǼ��[>�EҾ n�?���t�>0B�>���=�0��=3�a>��=(IO�#����4>x�K?@�5�(��=��#> ॾT�j>��>\�������Zo�>��>"���徯�b?I�P?s��>,{�>� ?!���������oU��&�C?5��21>=�|> �>��!P?�9?��B?��A?�Q?I�Y���b?�?-�۽pþ�/�?o��>KȽ���W%>�&�>�R?��*�l�X?B��>�&��v�=2翼t-<5�%?�*?�q?���6B���n=J!?W �=j�.?E>	�>�gR?� ?��>�{(=ؘ�?��=y��nV?Mܽd��>��J?T�8>6��$�(��_��g����=?=$��K�n1?��?y!.����zх?���>-������ݣ>;�=?T�+?����q4?i�w?l�=��=T�喿�׋?����R� ����u>t�>�ƾb)Ǿg���I�?�վ�� ��2?}��=#d���a�=e����47?�}L>u?)(x���F?��d�0p<�A ����׉z��q�!�������Ϳ�Yw�륿�0?����'˾0
��3޲=�c�>����Q����>*?�#C?`P0���Ǿ���=H�{>E?�>�팿�y�>�n�<��+�%z8�L����[۾�?�tK�)���D��-��>���E���Ŝ(��޺��ӝ>�,� ����v!�(w�>�Ǧ>򒋾�M���?���>��?]˿��s�������������>� �=]������q->�'?q�y�`���ᑾGA�>;h,?���{��>��9?�ᄾ����~Y>c:0�&8�>.�8?g�ҽqd=���6�������˾�,?� �dp�$�">�.�=b��Q����>
���;D׽ʨ>�L�>*Ai��{�@q5���'?S�־����Z>��=q��>O۽<�ɿ����d0;?����p�?�i�=V�2��tl�����Hx���J��DB��F�U1>�
?��:?��?����T?�C�<�y?a�<Q��B���X?�)�>�J��%R�{F]>��'`?=�#��+�?��4���k�A8<݈5?*���0���B>�����.?�C��V�}�c~;?������>®�>��;�]:9��0Ž?­>���>�=6>%a>�K��Yp��A����۾�
�
ɵ�ܑ?��b2�JÝ> �(>(U�=uU?��콺9Ӿ�W?��̽RžR���8�w��G.�J(վ��޾n�׾�z�?�Q"?S���mBm��V�?�Q>�>@����bg>�K?��@?7-~��@?o��>��"= �{����>���<򆜾�y� H�5�dJ]?sG��.�%>Y|Y>�՝=��!� ҉�������>�O)��i?���/?����L9>1�O�=n?Os��ﾼ����>�|�>3�8�V��d�>�?#=X�?��]�~��>����T�� ʾR�?6ӽ=��ʾz.��!�.>��?k�>�r>e��>$�7?�{�>�?*0�>Ř)?.��>�J?� ��?듽Ѝ(�Z?VD?��+=۲>m�x�'��(*��{�:���!?����5�>�X���)�YK�>��&?�G�AzӾq �Ώ��A�������3���3�+$h?AK?��=F��~}�>&[ ?���>�{�ȃ��	�>g��?��d�q�-?F�������r>3?�7��j�ڽu�S?���^�?�έ>ɾ~>���>\>�	�5b,=�8���
�V����_��0,?pd?��>��^�>Cm#?� &>�;D<P6�T6�>8]1?��.?,����6�?��e?��f��T�>j�n����>_�r��2��v>�>�HP��0��1?fK�>o/'>}���-���	��>-�	�K�>{����`�9?�(+<+���ؽ�V>)��>R	߾�;�x�3���?O���r���VY>o>���{��{C��X�ý���<�V��˕�ȩ�~�?J��C�9�2�=56�r��>��>�`>n�f�cI�i�>;�ս4ls�k���&>^;�> $?��[��5�>��?J��>&����8?r�=
��=~�O>J9���^?�
8?R�Z�AUs���?�z&?%�)>����lA��(c���>{�C>��!�?�w�E�5?�|���4��":��_>Y:þ��E�0�4g�>���P�^����=Ґ߾+�
������w?��W���C����=$�>~�?G��������C�׎�>l�0��<��^=1�j���?���B�?�g(�����8?���=]K"�+��o]�L��>��>�=^=l�4�j?Ӄ@?�w���0B�I��>S�=�g���=���<��?��"�n����m�>�^<��Y`�-h�>���>w?:YU���?�J@?�r澛��?x�?z�?�C��=�>��O�Z��>
��=�����D��>�N �ȶ6>��?!��>�R/��<�>����zJ?��t�%]q�����ֺ��v���9�Y}뾦P�����"*��j�>p��>�Æ�G�u�Q֡>I >�GN�����Y�[Е?-�#��VF��S�c�<;󒿿Q�=|C�>D��>
�����:���ξqU>.e�=��>i��>�4���i�v�/?��?7�2�~��?ɾ'�>h����>WQt?��Ծ��6�~�<�� ?��>��o�Ϧ��Ϸ����d?h��d>��<�	�>�폾�T�c���Ҽ>��T����ֺ�����D?>�7��-�� =&Xv�I������=��?��>�;>�Ǭ>,��>��0>�[�>|i6?��/>�t>�>=�Bw>[o�>� �>�#Y>>�>��>0۳=��=���P��9��M��ھ�Vo�"��An����ؾ��S?�� >]��>��>�d>;9!�[K��}����~>9�n��+^���!��-��͊>}��=(Žg��0>���=S%�>#�J��:���G���j�>P��&�Z��=C���r�K�(�⽣�l>��>��?\�?m�?��?��==���\Y����>C��>m�*��7m���>V�����=��X>�Ue=~j=0��>͍��yg`�hd�>��>�b>���=������_�� ��E�u�ޮ��8�;������B=�%8�����4�� ?�>�[{�=�갾�"?���=���<� C����=���>J�>�W<Y]-?��ͼ��>E@�I�Q?9,���3�,Y���?���>4(C���L�\ `=v�H�2oy�t��=���]@>W�*���F��%�>�@/=z3�!+\��$�����$�>/��&�d�=�N>�#�9�=���=vܾ�����c��y���rDL��v���N?`C�j#��6��nW>鳐>�/� )/��4�ڌ>���������>!ʯ=hɪ>Hh�[Gľ&�V�-T&>����b�=����Rľ�.F�0��>�匾ř
����>`��=&U$��8��۳=���=�OC��S:�c�>�tF<_�c>|��>޾�=��m>��>�[(?�I�>��Y=ES¾�M־��ξV�>�$�u�G�B�\=�_���X>Yz>�q�=���=�XC���7<�ϴ>) <ņ�&��[Y*� >�>�2>]�=�yY�E��>�*�=w��>W?H�f?lf>������=@�j�*���>��=�':���=��3��m�m�:$M����>+K¾
Ye�|%�>i���D>M�e��i?��C=C՛>QUy�������>2u>��=�F/�-zr>!В>[�'�>�P���u#��hF���v��/���>�ɍ��~�>Pdj>Y�A�=gDż��=&�>ڦV=�>U��> �3� oE>ZP?�>�%���!���>��=l0���K�>�{<>�o㾁����1�J����w��;m?T���X�=�D�=0�m>�h>pK���<��>N�����C�>�����⪽0�>���=�[�&��=��<?��>��g�DX>i/->�f=�0꽴���}��>}p�����F�uh>�=Z_.�nn��ǁ�>�>�p=������>w�>��G�}������瀾������v󋾴-��gx>V���ٜ�E�m��=�>u>�U�=H"@>�_�=�E?����>��>0�!�s�¾�xF�Zz�,�>�>�=y.u>���>���>RA�>��>t�t>�a?�i����\>��>�6�PI�>���>��?�����.V���X=��?V�8�]��>��=r�0>��"�i���;s>��>�6�ɂZ�o�xb�E`p>���>=7?�F?oh޾��?�>rx>g�`?�)�ަm��">�i�>-�?Q��>�8�BQ�C�b���B>D�x>�s�`�>���(���#�>��v���H�T��>�̦��;�>X�;>���lL��Yx>e}�>�[�>E>��5?D��$�=����L|��܁=���=T >5FѾ+J��`�"��]�x羒m��
��e�>}da�p>v��=���>�t�>IZ�=��=	�>�ʯ>%��<��`�3�w>��C>W|$>�;����>/��1��uH^>'��<����:��w����:��j����g���D>�A�=�	��30����> �0>�!�+�h>�:R������=
_>-����
?���>'��^�;�T�v���p>Ck̽��۾����>��(��r�;{>>C�Q���.��c���´=K %>8��>_�����=�E�>?/=���.9�>�J>f�1�c��Ե=�A�ؾ{�wC���A�g>�3?=��� ��hgi?H=�>�2�����>��)�'��iD�=I)�w��>��>_��>L��A!����)��ފ�>�\��ﶾ�ҟ������m�>��=O�h?�� ��D>�U�%�f?���z�>�^�:�j?|�7>(ҁ��g3��I�<�2>m��a���z:�ɭl>�G� [�Hu�BO�\y�><`�=����uS>G���J�<�_?=h^���X>OT9>�e�=!�o>��>={�>mF�<����=O�
d->iA7��j�g���g>�">����A�>�_?82"?V۟��+�<��>v!>I�뾼|���>�4y��3���:<�	�=�]�>�4=+½��>�_?B?��>���=�&����Z�>�P�9�����-=���w�̾���<Ω�-����>�H?t"�>[צ��츽����r'>�E���{�s�=4�u�!��Dn> q뼸�f�C@ս��e��2�>�ߪ>��?�7c�(�"�X���yS?���ֿW>�=�n>��o�����A��>,��>	�>) >{���=_����h�"��>��?}�����R>u�Y��)�Y�r��Až�x�>�Ue��E=0��mU����>�A#<��X��紾-�>?b_=N����!�=݊�=m�-��z�>���>
ɪ=.����6��^j���=r��Ǡ�=E� �ʃY?�=��Kh>�>-�>���ſ?Sk7>��j���>ݮ$?L7�>�;N��>g���Q@=�?%?���5>VX���\L=��i��(�<4Q�>��>���>�ah=c|پO��>&#����ͼq�=�6�y��R4>@-��xXO��Z8�"?=���{[����:>�jMW��^�>�cʾ��5��|M;�YW>�ͱ��`��~�{=_0�<����7�ܽ9(�>���>c�>}w�>s]�=NU,<�/�>=��>�^�=z]>���-L�:8�}������@�U	"�-��D�Ӿ8��>�u=����}��/�>
ϱ>��>~�;�E?������A=�:��K־��=(<>LNG�po>�+>Ay���3;�-�>��>�E)�j�ٽ���=y�d�	���=Z�>���G�̾�0)?�ھ͐� r?>���>�y��Y�f��û�d�R>��W����AX���>Ж?�aҽ�ɽN������,�pe�V�*��>S�^>�
�tg.���?~C�>F�,���p>�%�=2���lB������ŻW�o<!鞾�ν�o�>�۬>�s��px>���>=u>:��7}r=�f������=�FvQ�Vʞ��۾Y֔>��-��կ>~�L>��> >J��I���=ͿO?`e�� �\���U��펾���>�����0�<��=��>���-Ի�/�ɾ�;�>�M����=�R׽n?���>�ﳽZh�`
P?W�����5����=�!?¾;�T���-��>!W�������W�=�4�>�w�4�N�k�a���s�pK ?����#>N��� +�)�Z>�#�=t�H=��/>�����ۚ�r��>i�ʽ'[�>C�|���I<3Gv��W�>�&.��*��w�[����>QUN��)��M$L��1�>�t�>�0>3ko>���>�h?���>*��>f[�=�GO>�t��Q�����>�1�ӽR<,нׂ�>����;�/$?x��=�]�>j����E?��%>P8.�}�$��:>K5�YO0�Co�_ �==	�>�N��I����>�GA��׾���G�?%���:���?����>D;����,��wV6�~q>�����~��5k�eD7�N�0�ME�>V�P>4��>��+��G��>�/`>>+�=��?UH��=A4>����ܼ�>�5�>}�)���>~��5�_s�>+��� =B�<�c��\Ê�B_>}�佲�|?�td�̪>c�
�8�K=� �;�Y����=��P�ʾ��pjb���Ӿ�eĽIF�=nL� �?�S�-�X=e�>+�>уY>��4���>�$�?��?���>D��<��?)(f>�]:?�C�>o�?��J>��W?��>�{�:>%�@?��?��?��a<ct��%�>�ڤ�%�*�=�(��)�	��9 ?[�����G?��"?s6m� ��=���)��t�r�_}�h1վFь=�߽��+�����Ԗ�=p9W�L��=�<��>�7w�PJ?��@>jG��oh���3?���<�������F�T^�><���*�?�p?><(=?��?�
��ą��k�}��'?����
�Մ��6�?e=��-\3�!�0�'?���}O?�m�>������>�z~?twT?N�>6;�=*ނ����=��(�p�_�"�U\��|�!��?�S��9=��:��^�>�۽�����J��.�>.�h>.��s{���>��?��=m2�>N�?~�޽���#w=	1 ?�3v���پ����fP����>�XL�\��=�&?	'���-x>C��F�/�Qg�=z-��� ��C$��3)e=@"�>I���۱>񡯾�R�)��*��O���?T��.�o��+�tÌ��D�>�:#?at}����xcN>�Q?̱,�t���-�W��>���>�Bm�gO�>ϡ3���&?ƀ��)�>�)��^^?���>� S?h�>�tN��'��Z�>��) �w"B������=�s�\�Ki�>�5�����)�T�l�MBg�����A����=�V�>>��>�����>n��>j�]?��?�e�>k�u�sNv��f۾�&?mwx���쾂/Ͼ��>��b�K>׾_;��C�?pe2>H��
5�;�>���Xܚ�K,��i�,��>_*�>��J���~>�n�>�s>�6	>���>,�!=	V ��\?�kc>��?�i�<�;Q�*k���C���y��?��>#d;��U�>��!�7{^����9*?���<i`�=�2Ͼba�>�ݦ?&��<k|o�ՃR=O@�>+�>�_�a�>`�$>y�A��N��!L��2�S�4�=i׽Q#�>�?}�4\d�$'�<�?vk���Y��kT���?���횾���>F��>�%�����aD&�55;>9�i>��=4��������>O�>�V���>*=�aV=L+�=4��>9�?�?�L$��9��1�?e
-��aɾ��7?BH��7'?�A�[��>�=�>j}��<{o>�Y?0a��6꾜A�/�_>Xf?�0��aX=BG4�{�>>栾8�ͽ��=��0���Z����5?*�>���]�y>��?s��>�a>1�
>}wB��T3�M'!>`��=�I���?��T����<����q��ʞ��l�=.���xVI��=�k�?�F>�C���]�>�#�>v^�>�l�>�	F>�Kݾ5i8>��B>A��B?��X>~�>��H?�Rp?�{���?�M?��>�h?B���׾}?/ �>P��>G��R?KBp?2��>3�I��� >P4�reU?�!y����>��>���>��޾�B!�a`ƾr���?�<�%�> �A?z���Oj?_Z?u��<"N?���mn�>.�	>'�k=W;¾�0?&��=�U�=��>��?�:|=�A����>�=�� ��>a,�>ιB��B>Sդ�F���M?��>Oq?\pA>�<�?�"?�q�>�X�����>���>~4�?��X����B�7?9o}����in5����<�âͽ�τ������־��W���<�w���(�P!?�=>'#��r[>���:����o�ọ����>h���\{>Ւ��@s>|�d�����߹��v5?_�Ҿ�1 �C�����Һ��H	#�lT-�e�>W@�>���>Q:־�(s>�)D?��d>2K���>QR�>�F�>���q��=�2}>��>j�A?o�1�(�f��I$����?��D�Xll>�kj��X�?�N,��\��w?�:�?p$��R���������rI>��>A��Q-���(?Q,�>��?��5��X?F�?~F���'���B���־Ŭa�xN;��{>k�=W�?�N�� 5?�K?,�>�f��݉z>�e9>��?��뾡kf?�n?��t��<A?��mMM�y}�����>�=�ȃ�Q�=�ʂ>��4?X�	���ɾ����o?�\��Խ*�:���>��YwE��8�����>�(f�����b7��b6?O�=7{��k�b���*���j[�=F.���>��?�U�=>&��C�־�����O��)^�:�*���=e�������p�=0o�;'\>Xמ>?ꭾ�.b�����>�i�]޳�Y���>�.>'���n�>��!?�>�h�Y�	>��>�<1>kl����f~��Bt���_�L�Ǿ< ������=t{�AG�>;r�>|#d?SQ|?A�>�K>Va7?L��> �8?{�$/��P��>��:�2��� �e�jD=UӾĨ��i�ʽZ���^?�6?�?���֧?����\VE���>�>��l�8���錿��;�[�d?����>c��O?���>ͭz��	����
��?(�?(O^���?cz?mC>���BD#>��?A��>�&>��=V��=��b���/�CyH�� �dY�=��>�ھ蕫�o7��>�6$�ڕ;���>��>��b��P[�~y>�^3�ݺ�>3�J�?�"�>�)=�7>6 �>�ɂ>La�N�����?ߡ�>W�����d&(�Sb_�OV"?��<��{>|��>t��>��?Ф2?4Ev?��?���#?*��<���<���f?��9>5`>R��>r($?0ٹ=��޾���<�&�)f�����>*ɨ�=����y0?�WG?�J<X2��|Y��s��� �^�;��$�>�����p�j^οc��z4D?<��=9�K?{�����m?��e?L隽�`��ܽ	�>^�?�-���־`��>���=���>�d?��?0L�`B1?���?x;>?P.��*YA������l>@BĿ�a>MY9>��KrǾ��D�k
R?���>��?;�J��z?Љ�=�c�=�ܠ��9?1r�?\?})v�Qkt>��3?��h��E�N�'?�#?�%�q��þJ?l�"?�m��u�>�I6?l�=Gww�j�� ZԾ�ͽ�|L���>`�-?:�Iݾ���%�pO���+�.&�>�	;T,��,h���)?�P�=� S�V��>XSF�sW�S�վ(�;���l>����J%?�4f��т>��@>9�?T�D�b��=p0@>�}?�>������>)�>����y�>�Y ?�o>�
�� y?;.?�I�>�����>���=]�w�|<"�mk+����>��ȅ����-�+�5?W;S? ��>�v���[o��?]�0�ݸ��^�����؉t>l�>&2:�I:Ծ�N�E%񾮧��
A����r��=+m��ѓL�*<���g?�g��?�<��(i>;m�>3̰���ü�de��撾a@.�%�'�;[>�}������s���l��~?�
\=��꾎�>�h����x=ώ>��9�Vo�=�M��/楾A���K)6?p�8?-A�?���; ��5��ܵ�>��>qSP����rɾ���>�l��`I)��˾-z>0��>�O�>��!?�=%>�'<�P�<�.#?�P�>9����m =g�=�ګ�
��=�?i<@�_�e�ŧپ���<��>���G��ix�> \�>O�p�..�㻔�l���\ྫ��>!�>�޴>�H���0v������?�%\�C������W�>�x�����>#�
�߳?����O����<q��>p���k�(��{ﾫq:?l#�>���y>UW?������B���D�yk߾K�޽���>��*���(>ڭ�>�'�>�b���{�>�.W��;�V(�>'C$>g�>`뉾v�վ�+�Ui?[O����?l|���>�VӾLF)?C���$��*P�˸3?�o��Q��ƣ����¼\W��}�=Ϸ=�ݨ�����>[>������&=�๾���TNb��b����>��>e�?�K?P�*?�g>F7A=�R�>���=�B�>	[>`�Z>�t+>��>�m�=�Í>'�����> ?��>��2>¢�>`3 >.��=�SL?+)>ݼ�>k�?b�k;H��ƽ�{�8�̽g�)<��>aX�>y��=��;\ڃ����>�g�>��=Y�����=��<���w><���="j�>og�>�Ez��=yE�)�����>\��>zb
�B2�cn��X0?���=A�̽.Y��?���>�x:>�2�>.?4���>�.k>�!�>m^�=�j�cܲ��F�>�/���f$޼�,>$\���ց����>Dn���Ŷ>Os=�!�=W�i>u~x�q�>%� ?�����`��u�>a �������k?�-�>�̾�PY�dG��6X�����>�~u�p'�>~a0�jǸ�Z[1���>V�L=�V��?�f<�	E>'$������͛ ?�W۽� �6���=��>½(���;�J�J��?�>	n���L7>���;�7X���]Ч����������^���QҽϠ����L���>�0�=r޻��Zn� ��;��	�,��� ����Y��ߓ�Ն���<�-����$�+�>;��7�a ɾ�F?��"���=��9�@����򖾰�D>Wz<>E��b��S�:��s=��;��`?&;�>S��:j�"�l=k:>O ��nN��
jؽb0_>�=�>,r�'<m��!��t=E�<\�q�HL�ZM|>a�>~3쾽�>��A> "]�K�&>ՙ>��>�(��i�>Z��� ?��"�>,"�f�S��r�=��9�r֟���˾XMt�.$�=�T>�*��-�M=�N�����_�f<ZM9��1�����玾���>��O?	����>C��>�0>���>�ZS���۾L<ڽTz0����`R���P?�þ�^H���q=nj�=��G��>�L�>��н����/�>��<3)�~�w�=)�=��>�=��`<=�9�>&��>��T�b@�>uB���ܽ�ǉ��H�K��a*��Y������ˡ=��7�HA���	���Ƚ�&�L)>���>m�Ľp�>�y!��U�=$nV>�����?(j>����m��g?���=7�D?�w#����C�]>���W}n�����"x���o>[�>�8>��pJ>��>���gL��3�<��T=�
�>��?�E;�r�c?N g��n?5`�>�R��q4?�'��%~=R�ݽ��?B�ѾG�<N'�=Ґ��5�>K�<�[ ��4���	>-  >�S���<̧6�YYX=�^�=ҙw=���=�+X>��Z�.��t��9��쾠l��	o�=M�>��ξ�����A:=u-���R>`��>	-F��߾��¾�M��f�?9=Z>�2>0�$?l��=�ϾC��������?� I��P��@�>�v��t ?�Y�=0G����>��>�L�G'?h�<�_O>\��>r�F>��B���-�Df>A?�yƽ�K5?d�=��O<YS���aS?�6N���%����8>B*E>�纾�ì>pI���I>��>-��������>��>�=�Kp�n>y�?��?)���4zz�]�<�<?*�>c�=Ō^>e�!��!�>&�>UmѾ���=ּp��"��m�h?p �>�'>�̀��� >cV�=�a\����>S�?�$���?-���	->J@4<�V�?b����4?��Ic��_5��YG>-!>>��f���ξ��4H�������4��j���>I*�,��=#�r�\�D>"�p
`=�WK��-�>��)?�/��>Խ����1�>p�:>6s��>¾�$�{_�<�*��+'F=��z�����޾q;�>A,�=�:2�ĳ�	h����	>��>�X����'=��?h�>9���ʄ��2=���>��B>Ɯ��,�hN����==�ս�l��xҾ�>��5��ND=��/�Ni���#p���ɽM�߾E����>�>>�{�<�7xҾ�4?c@>D�龘�򾫇��2{\>?�?��<0b��x�繾���(d�>`g��!o�L�� 1)�;� ���>mї�=ˈ>�$>����I�!����=`��=���>�߃��?)��>CN3<�Ň;s�þ`�>h��><�e�����>"������CӍ>��y>��k���a���?�/�>S|���ȷ��	?�� =�>;�ʾ���>y<#����w���4\&���#�=�2�1�4�'�G�Ӽ�����/�dX�>9����������U��'���_<5�]>J(�>�{�>~l�<z�p����+$1?�/߽Q������x�=@�><�F��z|�!�>l,�7�!��q�N��>i0q���!�`뽾���� �-><����,�5>��R>[���l>d�� y�>�e��[�9��4�><89�31?מ�����3S����W>�uq?���=�x6�=Cý�SM���=�a�*�e=y.>�1?�	j=⛫��	>'n�O*?� �>0����j��"�$i�q?��-�=�/����i>y�&AL�4�>8�,?GٽK��> �V<���>;�I��ŗ?zl~=/Z�>�U�>���> ȉ�hi�;���#��O���Q="io�z�#�*�����>��I>zW��E���#?��ҽ�d�=Y����>�Cƽ��<�|��;�>�Ȗ�m���!�����>���>?C,��@����D>XB�>��(=�bϾ��>�;��=��R�p���\�R�G>8����"U�>F(?�i?>NN	?M�}>#�.>�ř>h��>�w�>}�D?4T=) �<��>���>[�>���<ҽ8}=�K�(馽{eֽ�S'��4?�:��!�_�V1�>�D��c=��>���@?%S�=w"��J8���y��þ��=�����W��9"�Z�U>`
�g��o�>�s?�~1�)f�>|����[�>����y ?����>��R?6��=B���=�v�Sn�>eI?Ŧ�BN>j��������<�>����	��=��=���Ν
?��
>�5�D��=5�ۆ=�
<�>tD�>}#�UM!>P�����>ˎ>>���?�7Լ�|?(��=k߶�*��=V�о)$������>O�Ľ��4����>g<�>�	p��5���æ>`v=��*�� �R�e�:����貽�u���>�ʗ��7 ���G>�s��6��:᪼R�=z�r����ď[���վ�<b�����d�۾�<�􊾒���4�"����8�Rҽ{7>b�L���>�as>&�>�Q����x>,
�\�ܾ&־���u
?�>>~
�b�<���>���>�<L�&��?���>T&�wϹ�/���\b?�`�>(��< ����n�=��D?��T�����P��=v)?7K��!>�u��Ev�<!�I2���=�l���j=ڊ�=��¾Z��IM=����\�̼�=������w�^�����%�루�����?��y�y�����3>8C��B��u���-��v�;����l��=�F������U_���E�<?7н��
�>�[>U�޽�pľvf�4�&>�pZ��<)����Md`>����������=��>�a��<>���|}���>:=��i�7i��j�}��p��)�>I���P�>2ﾃhm���o>p�o=>�a>C)?D}�>?�P ?�Q߽�R�=�"?��D�^q?*B|>�[�>PFR�E�ҽ�����������r�>���>Ȕ8?xĻ=W׾͗=�T՗>�+x>���=���y{���YQ��0��4��>�vཉ���R��a.l=�W0>�����F�5�=�mǾcJ;�J荾��Y���4�}��<`O,���>�,Q)> �>�Wi�f�?�JA��U����?��>gO��O���{�+��y��m�)�>zj�>�����Jʽ[].>W�=�i*�N��0
+>֓�=����+>��`;���>����9*>�����,�"��>�.Ӿɿ$?<-?O�^>�����I>O(��l�=�$�>]�Q�����?c- >$ւ��!�2�νW$?ʓ?Hno>#��>La��34>��|?��N?�^)?+��>��H?��}�J��=,e}>[�!?w�>]C�>w��>؟L�n�j����>,)�?�����>`?�,>ڴ�
�������?�R�7�j��>'nJ=^����?T�"?�ߩ����n�>���C�>0轷��~�?n�>\x����.�>���=�LL�w��?8eP�$�6�g���!?`��=s/����ӽSL?�^��Ur�<D�ʾ��9?D	?��>�q��08?�m8?o��>�Y���o?����Z�>�����vp>��>��<�3|>�f>�"�2?���<�����u �
��>?��?�\>"�T>3k?WfM?���bT���v��j�=���&�J?���KmD=��>��*>Z�ٽ�B6�����ɀ�=Xh����#��B�>G�?�
]?�s?����7t?�9�4���H�8��?���>9�>��;��f>`־h�gi��0;?��r=�c�>� n���j�Ŀ`?A�=�v�0��\(@�Q�=�*��c!۾/��p ��(�^=3��U������t��� ?�	���>S�>6��>�ɾ��=���0��=%��Lꎾ8(���7;?:֒>�A)�*�"�������?P�о��8�R
�y�~>$��?4�w>���=�l8?�``>�;�>R���_p1��"��NI1�u@?>k��:��%�?��3>y��N8��!?�>b#�=L����֣:r�>�@��I�뾽���;>:6�;k�)>��E?:�e?8�>���������{נ=��q����o��>~f���Ҿ��
���^?�$D�dТ���?��>��_�#�V�JPf>�q1>�2�_�!�=y?!.>[�=Z ?�T?��E��þ���?I��0���<�>q?��$�l>�]¾������?脽�\�>D�L��L���y��?��s{J��Й�()����'�<n?�g>��>@�~�6] ?�r�.%��2ً���?�7ֽ���=㎿�䤾����6:���v��?��R>>ؾ[ݾJh?�1m��G�8�����)?�GS���E?���?�Ơ�Ә�=m?�?""ǿ��4��b�>0��<� ��9�>�x�>����Y���G�>޹7��y_�1J�?e|h���������Ba?k�|>ErϾ&��>���?QC;>��9>���>��?�Wc�O_�=q��>y����?�>L�F?�9�?��B�-ڽ���l?�y�>�� ��Ԕ>�:R=Л�>O#'�H�{�*�?ò�<�=��|����>�]�>��|��u�>���<E=>)��<�4
��0U���<�I�־Y3�?h��N�þh�?�9�>����0��E:�>��E>X�`��i&�|�?w��>��>J]G> %?DQ���=�|�>�Ȕ�ٶ�=3�0���?V}�?���=ɋX�u%�=o�s?��Y�r<�?��?�C_�!w[>�Tp�)׊���x�8�->1�D�Թ�>��V>$je=;�Z=�K?��:�:>=G�����>Z��>l`��7?>5��o��fQ���*^>�)6?�]L?�	�>,=R>�^&?yt?�Kf<>�A��];?1�W��D7?F��}�$���,�p���.*?�^=?��?p8�=�'?5>?I$����=c3ǾO�?ȃ�$�>y�+�0It>;�<�l?.&���=E���o��%�>�>���>8�>���>U&?�־��>h*7>'1?�����ξ߻T?��?K��+k����Q�z�Y>X���,�>�:�����D�s%e?���l¿���f�>oO�?W��a:v>Mr?�i�>I/-�F���..	��b6��4��b���Ƚ���>DCP�&8������>QMɾTV=���I>	>jg�����Tvq����=p��>VL{>��>�MK>!G?S��>��/�*�ɿP+�>�(	�� <�~3����<��7��6?�8��ľ>�����БV�:���_�'�½Z,�?0�*�Ht>A� ��?TF�eB@>� �>B�?�iS����46�8	�>��/�C$6�[���3�>\�E�Ǳ�>����ѷ�h����F��@���䛾��w�U�>d)����sd�}?��?Nc5>��\��WO�.�þ�9���x��cu>\�s�)	=ʾ��$?��Ӿ��i>��W>ᡟ>�j+?�|�>����H�p=��ɽ�c�>���0(U?[0��`�>���GQy>�TH�y|#����	��)>1�o>��>�߼M��=�j�=I�m�ؐ�h�|=O���/Զ�F�O?C�6?��&�� ?��@?�i׾�����3?WI�=r�� ��u$?�Ғ�ӊ
>r?�[S�>�?碒��G>��?��>Xw�M�<W+�=�(�b�>9�CM���T�>]�>qގ�r����>�K ?x�=���?��a�ͽ6�ZWU?fn���2?�@�>s�z?[G>l�E��+��?����ھ��K?5�C?y�����f7�=|��?,5B>ۦG?��>��?V|��N>���#�󮰾��ܾ�޾��^�X�7��ch>���5��=�R��.��=�CT����v�_?ۜ2��E�=���?V�?����g�Bŧ?�y����#>��>�k�>�̔<�l��?>��=Z�S�oO?d	?���>_�?�����ҾǄ?+�=#����mJ?c9?V�O��T����=�WP=�J>Ic��}{�>e?������=:�p?@�<^f�;H�t��O��ġ���뾇��=X����&�>�y�>]�?39?1^/�8��>D��>�F{�]�?{�\?��>���ƣ��<:�=���[>4ȴ>��=��>(�q>}����0?g{*�G�Ŀ{�I�lC?�� ���\>2��>��p?��x����u{.>�6�=��G�I�>0��=6J���?d��� ��Y���x�>��<�ʛ�srq��\?�7��t���N	���J?Xy6>�2?��U>8��?��f��>�*�?dLc��tR���B?h�-?Ɇ�>�G>*q�� ].>2���۾g�R>����>�*þ�G?p =��ͼ5��q����Ml>�O?��ҾI�?�M�>�8�>Õy�6��>(�>�D��|=qK�>O[�>�r������)�>x�q?�K�<�1�2�
?�=�>|����>"�t�,0b>���=�J#?��a�l(>��=�=hZG>r�����t��-K?	|�e����G����<G�>jK��;���֤�A����C>m�-�󩼫������+B >�e�[=�H>�y:>�Od���$>K\�?�û�*j�@��>/nC?󯵿�����>iE ?qz�lp�=���>5�@?�XW�(@�{7>�M�>l)7�ķ��j2�~*Ἠb?�$���'�>�t�>h��>qh����^J�e�����>��3��X�=5����.?��T��������.�>Eٽ=F����о�M%?F�������Tn�=z�'���]>\�_>�N?�)V��n>c�H=��=�v�=s�3�ƍ*���?G��?.%�k@5����Se����r�?�y>A��=�:�y�?�������=+E��>���>��?�@?��?�+?.$�r�1>�2�=�b?��ɾSM��>��>�F?V���>��'�޾Y��=�e�>�������<o�X>���>��?�j?��W�?
�>��>��f�Ċ?k�j?�Te�/��=>�_?�2꾃�ɾs�1��ֆ>���>��?
V8��['9��4?��S>z�<Y����>D�>%���5��>?i龝Bξ,��I\u?/i����>9��=����b���>��׽8����$> �����L�bI?��(��������� >O���߁�����0e����ӱ?ZA����>z��:����ϴ��Mr�3G6?��8?�a��ʳ���ʾ�\�>��>?WP�>�!��������7��v��}�����La�Ρ�~[��	���7�7_�X�YῼTSr�,�a�"cȼ��m�����fc��e-������B���u��ý HQ��-�;J�=���<�X�=�����<l{=$+�<���<̀=�<P=�3=�l=_&d;3V=�4(=�Z�<�D@=���о����;�~=��j=>��;�&�|{g<N으_[����<�7��i�<]���N_���S]=��9�N=��$�nbs�)�~�I=qJ��3ּ]67��=��:=������G��w=���:Z��;Yr=)1 =Sf��¬���f:I��=�>3�,��h\<��.=�̼�M}��fҼ�O)=���<Ԙ�=��`=:F�<���\x�� �<;�=�м)ૺ��2֍<<%n=�P�<($�<vbC<��< ��;�=��VR:��=(��<v����E=-=N<v�<Y���8�������Kw��@���j<@�o�����@;�Rɻ���F����ػ�����<���<�c��xS&��<��΅��(^j<�o���G�Uk7=�s
������H�����-6�<	^��Ə?�ԓi<��=���<r���H���/�:~�G��p�A���!=p��<K;�Y�u�,�=�e}�i�p����⚼a�w�ڵ�K����~;�/�����D���?;v���m'���J���C@�<6¼�䴻vc�Qzh�V)�<ed��S�=�Nݧ�x:`�Ϟs��F�;��;�oR=E*�a#����s��<�y�I���?l���F�t�d�Dj�k<�<�U8���i=7��<�Aۼ�Nϼ�$=�M�;V�=���c��= �	=��{< u	�{�*=���<�8�<���=Z�<��弹��;>�IЄ�R��Z�)�d�W%a<��4<�zX��\�<?9���-!�,�(=9#�U��=-�[�=�<�"���)���|�y<���<�BK=Ţ=�9=�t=?��=�����e=����������)����ܳ,�P����<١���܌;ʂ��|=��eN<��<����Н�~-w=��=�.h<ɱ�<?�#=��=G�޻l�b��I=�򼍷�<=+�����=,��2��^�:���&=z�1���ʼ�7>=B=�2O=D*x�˚<)��<�,X<ZR���<�ܳ<9�W<�T�<翼�L�<3<9�7j=�蠼���<����(.V=B��������#��vT�K"a����<�s��6f��^=��W=��$=�e�	�^-����u=!�ؼ��D��s�� = n�=Gd�=j�s=$j?=e��<�e���]�� g��5H<8�ļV�c=�����P�<�K��1�=�ɒ�"Ã����;�H>;V����t<pЎ��}�<�.���=ӺR=�z)=A���=?���=z����_�4;/�"����]�#��p�<�	=Kx�<C�J�ڱ!��[��X�G="��b��iv��(`�<r�=�2)=�-1�Q�3=5n�<~ⅼ����&�T�F=D�w=2���9�<�P1:��<�Ym=4�����=�n]<���<ې�<�뼉���y��=\�<�/���|<q#'=��6=�mS�_�ռ�nK=P?<��m�F�==��i<�yN=b�)=U�]�9������]C�;�.=�m=LQ�<�]�<g�J<13=C�S�'��<�̩<�`�<m�N;\[V=�1=�(=w�=�c�o�@=��2��n?=���ܻ� \=�='h6�����/�������<Ԉ�۷�<^=O
9=���q;�H+�W�D�G\;��I�;��_<�lԻ@��<V���@�R=�G��*=���1Q:��%#�w(��;�����9��R<�<GI�f�ػ���=�ur=I��<BX=g��<�3�_�_�H�3�|EQ;G=$!=�R<pc=D0��h���#�׎Ǽ��$�9�/��i���cy"�B��k��=�e@<a�<�&�7(u=61���0��79�9�+��Y��ס�<�G�yP�Zm=:�d�L�n=-J����U�H� �6=eθ��%K�8W=�Z�=Iy@�9�=�V�9��0=E���g���Ȍ�\���b=s<}KM=+����u�T@�<]��<��j�(���,=-]�=,��c�;�#���1��E��9��/�<<m�=�h�N��{�}=�?:;{R�<�����6 ��}�<rF<���PBV<j����$<<]s�+��<��k<������w�)=�B,��Q�/��"0���]��s��|�ν�d6=�~�=v�u��N<�z)=�e���/����ž�=;�~=i&!������;=w9*<�����<��[��������er߼��=��y}�����g�$������\�;�L�M܁�6�� ���zJ��R�χ=; =D#�<��;=I<=Q�м�۫<�z��;܈=%D
=D܃=�Ù<g�(=�)�<�E�.�==2�'��<�6�\�O�� vp<jU��v�J=*À�-/<�,	�e�`��ǽ=��<�$��4��<W ����=Vm���߼�Kl=��p=3�]���<�9O��>=�3-��K�;�耻*=:�P=�*��~=���͝�<��U<t4B<�o�w==C�ջRzJ���b�&�*��I������G���x���h5=��=6H�=Y�6��;S=��<���<�S���<��t<�U=нP<L�;�߭�#�Y=�P���?=�ٻ��m;	Z��<Ѽ�-]���o�+o����<�b��>0;�J���[�H�,��th�9@a<�Q!=���;e�<+��(�<�T����<P�K<N��<��� a<�N2=��k<1��;@AW=`8�<AY�#�<�M=��<�)��Y���e�;qI�=%�=t���a�<�R=�|=	a�:�;z=xAt�/,��)�<s��q:��;ž<+��:1�=OT;�WK=J�="��<��ȼ�ԺJK�<_i�<G!��:<K+�N==�C<e�S�����L�=�f������E�_L�;Ǐm;���G%���+�I]=��=н=G���ȒJ<��<��&=��(�.�<��;-��=U ��<��;B�=͋�<G�ѺO�=�|��G�$=�m��&�=�4=�Fo����	8:=�.��M;ޯ��+�����<��r�l��<�ɪ�P�^=
m�<|	`=/���q=<�>��}|�;j<,�X<��Z=��>=+]Sk=�j�<������ʩ:LC��p=��=(40=��"���9y��d&k=����s";������V�ϡ����C�>e"<�l��b���|�*��<���V�u.3��a�;�+q�ްf�T�F{� ]+��ꋽ�����B�7j��Oo�턍�h��;c���2�:A#�<܀��F������Y�B:=ۖ����>��J<A�m;�
'<� �1�=2�p���K= l���%�</"�=�=#�����Q�h��(3���7��n�M�3eC=�fq=��Y��ȫ�?�=Иu<x:�<�[�=k;��D=Z�;��Z����A�%��;�=�;���<Md2;�>���.����C}�تٺ�m�>��=�̉�b��,5P�<�<��;����׼s�<bԇ�F�,����q��b�"�o���;h����<, ���������cS��t�M�C��#<�����oK=�k���A�*��:�hw<����Q�<�I=� `=���=7���n�<�H=�|K=(�%���p�%�ȼ_ <R0=�+̼l��;��=�&�;V����Ľ���F]1=�� �ޛ�<�Q=��=uc�<ƫ�<\��<�"�?Je=�0���<&5�°
��gr=��4=�f��M-=�\�<�=�2��xw��Ɗc�qt5=�.i���w�7^ ����<��������JE�Mc3=;f9<������N�W��;�W�<u���R(̼�b-������J
�� ܽU͊�͘=�1�����:$�f����,��U�L�������� u��ޢT��	�;J�<�(����<�W2=�x���*5�a�X�h�<�I�=�Щ<\��b)�ˈU����<��<��Ҽ�nA��,�<i��k7����v�dl�<_�Z�f�{��B�<�|t�؝\>1��<І��c�>	VD?�ѧ���龿4�=�߭>�T�1����"ս>Z�����b=Y�>)U�?��?�`>f�>?Y�?�U�>ȳ���<�ag?u��>^�	��s���?��)>��,?O�⾣��>{'�?Tڽ��a>��>�wg�x��=?U��֠�tb?��>�#8��*��᯾Y�?�񴅿d��>_��]4?_+�>��>|Z�C�:�`>�#�>����;���K3���t>�j����H����>�H��i�?�D<1Kӽ������>�m?�B?O�e>�"�Ŀ�;���>(�����">��x>H�?Y�o?�>S?��?6�>N���&ɾU�?����>�m�>0�=�����:��>��>=�����;�>�,?Y�1?-�>�
��.F�vl�=��?��Y>�.>�Y?��>{��Cꚿ8�ƾ�/����Bu���ӿ\Ⱦv������?�F3��<Y��O��e��>�<��Z��E��(�?����}>��?";�?��ǿ���>vY=�߃?���.m�����	`�? �п�����
.����>�r�������ǽ�a�>�M�Q����4P�,�:��a?�kھfԧ�¯M����>�h�>�'�V����<�3��t3���ʰ�'ʳ�����=]�M?��I����xn%>��a��|~���&�L& ?�O���m ���=��;�kf�>�	����v��r!?�jL>X�>����{\�=��>U����FO����/2I>���kYZ�lࡾ�6?>JB�>��>}��c <�up=9��>���K;��W\)�R��>��$�3T?�(?tn��='?O	�>�h>
̵�;���>���������ˉq�e6?x2����<~���1����4���~u�N�]?B�X?��%��}2�2���̊�=TԶ>���=�Ҥ�>Ko$?/-�>��'?w�?m���{r?=Į� ��>a��>��ľ� :>mmY�´�>�<>�v���5 ��!2�cѾ$:����
?��i�Z�>wS�>G��~���4�?��?�{>7Å�>!�?��>u
?eV���B�>}�<�fi�<m�v�����K%Ѿ��C<K�X���<}�?s������v(>�����?>�S��>a���,>}�?�C��
�r���Xwy>� �=���>�A[�pf��n>�>F�>qm���%�h6�>{�̾���{�����c?0/>�#����zS�a@�=�G��(����[����>�B�>g�`>�Ѷ��x�?N�B?��Q?�T�=�����]?��;>[@?�� �Z����M?F-�>N8�ը�\���-��྄�>>��)?@U������f���Z?�z?��ξmI�<�Bf?MP�>�G徱���.&�>m^&��˟����<��L���y?�~?�Sq��̾���KU=
��>0��S�j�|?�S?�q�>�c?�_�?���v���H�n$�J���K?���!}$���>'�A>��D��ľŕ�>�����&U�a�Ⱦd8�-GW>y�>��c���7�?�3c?����0�Y%?j>>�Ȗ���H����?������嬅���0���U��i>�>�/�<L�>����^+�7y�>/�й�<���,�=-$/>���
�?�OB�t/�>�`�>ަ��??�T=f8�>c�]?��%��H�?���<=U���$���j??��=�ž:�=��
>O���S��.8�?���>�v�R���&;��B�n~����#�+`�?)Lb��٦=O�=@��Ci>�"L=�g�>/ھ6�2��5�)�?�3���:���7�6��>�7E���)?R�?�L!?�'f�T>g����>t?б�>�gx���=�l�s�>qk?��>j(�^:��������*=�"�GV�}����v��@!�>h;?J��>3���O���>��?ĸ��a�>�8?�u㼹 7�?þ|>伜L>g�׾���w� �*_޽�ې�2Y���H����о\�I��_'� �ϻJ����3�Ɋ���>���>
�x>�<m?]I�>�F:?�'M�rJ�=K��H��>�+��f��b��>t)�>���?QS5���|�Ӻ꾇�߾y��=���>�=�\Ⱦ����[?��=�6��6삾[�R?W�}=[6�wX�?��]>A�?`w����̿��>z��}�����"?#,����>3����
�<3�ʾϡo�=ȁ�L�?ˀ��f#������D�?;�n���w��Ҿ���?�R���>N(��]!?��g�ɓ۾�"��OG�#�A�W_�=97��]8T�酌>�W�����h�Pz5;����fj��$���p��#VӾ��3�G#�>
��j�K?�h?�*�3�8��a�g�>7�>�ݩ��A��?���=�8�����>��>�*�=��پ�1=Fe=�+?,�K�	QN�n�>�~>����XD�I���R=����҈>z�>
%��@N�f=,�]?8�#?�H�<	�7?`̹�\��>,-�;����������?2�{����>4�?���s�>0^��\�a�8g?v��`��=�?�?D��Q
?\�#?�1 �t]��O�#�#>7�Ѿ+6�<�_�>�]���e���^�?@��?���>]�,�-j�?9U�>`�?i���� @���?��N?�ă�����w?������=aUz>��c?��.?7!Q?������ʮu>��޾�(�����>50�?�S⽋S��#P>'�>?�#�Ce��F���٫>�?�E,�a���&�K>e�>;�5���*?���>TV���w��K�	À�%��"�6����u[!��^�=x��&�E�oMG���l?q�>Ex�>��q>G*?�t����/?P��=��V��i=����|�>dܓ�X�>{?r%]>�Qt?KK>T
�>ےy�wH?7�_=��?�E�������>0�E��?�4�Q>)���N6���z,�g{R���=��B��x뻇��� Y�>|B?W���D=�(�>�?��L?.�!>nϽK�	>��:>�b��h>)��<3�i>�����?L+>�`F?��p?X��Yf>�6���{?P��<A���������G�7��c?Х=����<�m��ݼ������}?ֳ?<]о%���
�>~�x��a���\����?�� <�J=�4�>�x�>�Ⱦ"ƾ1���?Q�$?U%u����Z4>�8�>k�>�9��>~�#>v��'V�>t8=X�ƽ�
v>�4$?`m�����>@�6>�6���\�|$�>���=+�߿A��>mB>8�b����y��j��#ѭ��Rh>�I�>tt��K��?��� �ؾl���{?�$��FJ�z���
��=/�9��]��d��>D&>�Z�>v?n�z/���i>�w�=�[X>G�2�!rO?�6q�Ȇ���PM��N-?&?+��>�{"���?�?|+3?�ۖ��gu?w�>o�J?ʂ��$#?�v�?4�&?��$?X����H�����=&m�>�����J𾏩}>���=@f�>$۝=v'?@ ?pؿ|���=���Ř4?�"e�S��Y�>�@*?��������>��m>��W�b'�wAU��[�<f��
==���:m�R=X>��>�S�>�!�=<}�����<n#�>y~G�	�>�D'���>,�;��ǁ��4>t�?r�?�n��C��>���=��	�|ۥ����|�H�h�L?PP�������٤�8e>���|��>�?�u�?�}�>��<>n݋>?F�>sjM�9����J&������7�>�?�>�H]=IΓ>F�C� ����ھk�@5�9?��?	}u?y�?�+?�پ�!�><�>�=�� ?�i`=jb�>������b&>�q���0�>+���[��>��@�-��`�h�2'Ǿ5H="��,	�m=
�=�>����x/�g����3���>�d�>+n?�ݽw��>��E>���>vv,>�<��c7?�~�>S��>x-T?D�$?� n>	�>~Q?��4��u�F�$�Y�=��?_����\�=�Bl���7?:��z���.=ٻپ��>z�z?��=��>'o?��ھR��>L⋻
�N���H�f=��������h;�i�����k�䄥>HF`?V�?��\<T�?� �?c��?Eg?�YE?ـY?G�%?O��>���>_��>6\?��>�0�?��>>?w��?��?
��>=���Kx_�ݠ|?�L?�/�`1>������V�������
|�<��=?�C	?~\�>��=�O߾�;>[!?�񂿯�7>�7��u���� �i�����"?o��@�B�����>I�ܾ9�O���&Y?;�ﾭ��p��>�>�=g]��>h"?���=9��= � ?]�?�gl?KuJ�?=F.潖�D?�ӫ>m��=�H�>r��>ԕ�=�ȾÃ����>@�>ta��Mt�>�q��-ǽ�)db>��>+��踩����>���>�"��J������-��^�*�E:��G���2-�=1�������*��B���>�hѾk���m3�Ƃ�}?�1�=_��>�L>�c?���!�;���mS?UBm=�RP��<���P>ܯ��e������D� >�^S>�of�,���^������{�:�5�B� �>ߎ�=�Q�Y��@}��je�ђ�|��V�ľ���=9M_�}o;�g��>\?=t>�觾��>��<-*='�8{Ҿ��R��⦾����j�@�@��@p�@D	�n��kǁ�G�=��뽳g��RȌ>���>u�F>��=��?�đ��̾�������*���	㾬��=܂�>Xr�>��>�>�νY(��RP�(��=��#�ƾ5޾�?�t*����r{?��#��P�>�1}����>}$N?��z�Z�
>Tm>P�=Ί����
�ݺ�x��>��1�s׋��?k>���=c?->_$���~�>,Y>�¾J��4 �ֽ�������g����U>��;?���IE�=�6:?�1?n�̾�/1;;��=�b4>wL��}T�~�M�ե�<,a̾o����#�W�����M��И�='@e>m���&��w�?���U	�B�/?��<=�� ?�{�?
Z);;?������|�גw>�?X?�s4>��^��˦�2���a:��`��؄���6*<�W��������*�:���Xy�=�O��\>3d�=b�%?���=�b��D��>���>�:?�]���>?��>��ν�m�>��պ�$�o4C>�36�Ta>E�t�>4��=g|A����`���L�>�X">4���=$>x�?᩽>X�>��=�?�����Z��:�e$�U�>�IU���?̒���۾*�?�0佁��#��1]��n���^w=�Փ=�H��8H>q�_�.Xq�'��>��>�}����>�>��=-�>�;F�n�V>�X�>��J�@�����&�=�;��圾�0���^���*>&y��2�g�> S1>C�?���>�e�>\c;?"�>��`���>���V��w	?��>�9>�.�?�4�?�K�>A(3?�Y?pa�?K�]?+Y�>�O�=��+�͂���	�>�~˾]~�>������B>H����O�?n8��V?��Ⱦ;i�?���?ʆ�<E�*?l}u�0��6Z��X�?�w>H�)?-�p�I�R=aS?4�"?{pS>=u�~vp?4w�>�Y?���?�s�L ��Aw>�U����8>�d�,�?@ �?p�D�oo쾣L��2�t�����p<?l�>�]�X6��Ke�/ >#�U���?7�1��>��ֽu6?"�4>A4�>�E���?��]?�ξ��?��M>R/�>�~㾭�d>fi�rd������pp�>_�����J��N	�A�>�:���ԾLs�=��ͽ�0�>4
=��T���=g[�>G�=X/`�����ȾǑ=�T����LF�`	�bq��m>�A�-�c�!�X�x���D�=����˩����?�c�@ �>Q��>�S�>�>>>����e2Q���c<�LU>O��,���,`>^:;.����2(��:>i����>���>FYG?|s�>r�M�����!��ů=R���.>X��}�>��?��Dl�� ��+��=���ㆽ��5=M�Ծ����(S�[���yھ���=�8��-d4�8�<>�z̽?�>��4>,k������B��>lC��*.�>�?��?>`l��x~���N?����&�>��1� �?�m���>��ƚ?��;��>iv(?ʶ�>!��=��?}r۾��)�lC��I:�͂������U���}?"w^��q2��(����>t�����ɽ����5�8�P#Ҽh�߾q�>l��=���=	2B������>�i٣�,�ھ�L��g�>��'>�s�>hP,?���;G!��j�5eg>��>t�_��r�>�?>m9��a���9\�B&?��c>N� ?�Ȟ>'����{�>t���lpl�b�#�&������$�>j7?����V/�ix>T��=xm?�z�=]��<��N>��o>�7>�?��H=��t>Q�,=��=�>r�dB���nS��Q��9?�,�>�f5?�_`�q���
?�U��>�<5�~>�K>W��>�!��T͠���Ѿuz�<�"��l�>��t�=����>�9Ǿώ�>�`>�AG?*���eE?J�4?�t?;E����?s}�?���>��V?�BL��� �����4�熜<J?	�>�"��O�(��b�������Y��Tr���>��>V8�>v� ���>x��>�|>�n�7���
R����>�!��
�w�>RTL>��8�୤��B%?0 �=ԗ���>5�����T}�>��ھ�q�>R�_?���ҳ��F�)=�?�"X?�s�>����5��e̼��.?*�?1�?5{z>�����ž^ǘ>���<?o�>xb�?�ܥ>��@=
cF��_?ϯ�>���>׶��z��|5>-��=v *�n[�\o�=�Z@=*[>�k5�p��G������5쎿��$����������^>II�.�Y?�<D?����,��>�c�>��g>�Gd��K?�)?z�G?f�Q��ݶ>֜#?xV�<^c?v��>᩿>��*?ƴ�=�L+?�V������4x���м�� �9���J�/���+�{���<[1���>��Լ$4k>OF�އ?ׄ-<�?�}(�X/�?��"?^���d�<Md������쾍+Y��[�>�Ǥ>M�?�,�=c�?��>\I��f�Y�6{m?�	?K�پ`��>u�u?R ?�xH:<�?��0�¹�=��H� 됾ŗw�.�.���J���>XF޿$T�?Zc=���)������b�۾a��>����)�>L�m��l��Nj�=aE4����>|���O�J?���>��Fr����>d,��m������=9d?�A��fl���?!���zo��?�/?uYx=�D׾�2�����8~R?���>�C>ܡ9>.i?�
�>�
�7�"?ș?��>���Ϋ>��>p��>��E?P-?ף�>�B�<NQ?\ʾ�0*>�7��9=��~/��p�/ZH��Bڿ?0%�M:�>���>��f?��>�C���>�����r�>��)�<N@?Tn�B�7�gW��9>G����U��v�a�h�L���=T�dM!�gY:����>yY�aGK�CDY�吉>m��>���)��<F���'.?,?E<5�֐���ξ��j�Gk���c羶���8?�3���s����ᾪ�?����˾��ڼ��>h��?4�e>�n�?��a?��=�[�"z���ã�U���u�=��>��>��-�ҽ<��͛�IsU?��?u|R?���>�x?�#?h��=�	\�pǽ�����>!^�k8�>s�˿�Z��F��3L%>mX�?�=��m=���>L��x�>k۾�=���:�оl�}3?,���G���s 1=��=�T0�Ь�0	6�9�����辨p5?ܫ�T�>���> ��>Ъ��=uA�>:��>��B?�J���X$�>Q��>(W����=�n�����>;�����>�E�>�k?�k���;�+�>�
ž���>�0�>ג >$���_Y>Ri���>�Nݽ�ݽ/ق=#d/���5����>�����/��(=�O�:;�p�g��>a�/?{cN>����y� ?�A1>:��>�-4?8�J?v�^��A�> ˆ=��>7�p<����?��>>���>���vؼ>R�>��)���>@�?+�>�2?���p���bW��]��,��>S�?}�2?$ �>�ۋ>��M��>��>�Yľ�z��M�ܽȘ��[C>�@v=J9��C�>ۻ�Z�?N&�>fq �gp�D�>�^!?�����-�SJ=T�Ӿ��m���Ǿ��{>>?�!�>yE�>��%?T0?N�q>�d�YB?�?�j���ƾ���=d�a���n>������u�b=NO>%�>X��<�V1>�e�~�>i>jQ>&|c>T=? ��>.�ּ:����|P�|��� ��B���u�gU��;���0?!�R=r�v=\�)�@H�>�Gھ�2�k5I���.>3��>$�>�OY>xz?軭<nu�=��A$�?	�.>yB���Ҿ�h>31�p>g���	��q[?�)#??���4IR>�ր>)�=*N�0��.�/�F��=0�,�2z�b�$?B�?��1�`����¾8Y�䬌��|����>��9�0#��[$��6�>�I�=k,r>M�S��n�>U�_�� ׾ZK���19?^=��� 4�]՝�q�V��@?��e�������*>��>�?��?��f?HW�W�̾R�^��
(�w�N���>p{�>��?w�>4�>+ Ѿ4^�>	o9>�Ͽ����
U|�q⻾��E>��I>�q���u�>���>��o=�	?�!%?���=^!�����=���>��a�j
t>,ni���p<U�><�N�X�q��Ee�4�`>Z�����=8������=���=K���ʰ���!;�����[��!{>Da>X?�\�<��?Y�7>�OJ?2��=��0�"I?љ�>��>/^�>4�ǽ�Ĵ���i���r���Q��1�=h.y���n?�����aʾ\�>x�V?'�P��U��Z��>?(�8�62�>b�>9�?�i���߾�>?�u�<��L=��	����P0�<�Q0�@�,?�M��2A\=;�>- �u���$q���Ŀ
�"��̥>�w3?Γ�%����1.�sx��y��>�e)?�Ol��c��S�$?��y?�����ˋ����>y]��)E������>Z*g>?V-?��>*�+����>� #?�脿@��l}�>�N?1��0�>wъ?#'D?*$��Zs>�yɽkj��'L1>�>�Ž��q>�\=?Ơ�=7�?w��=3h��(>4?�Cm��ޔ����ӽ��t^�7��>�1��~���>� ?��X>l���0�p�1�y��=$�z���>;����=D�o���w>�ͼd��]!-�:U��Q/��Kf�7<ʽނm>�4?�?)J.?P���L�S�᳾̉پkH�>XO?+g˽g|��W�����=#�
?+&Y�6�W>m��>�T?)��G�G����>�-?\ȣ>%#l��x=�DȾG��?��k�&��L� ?:�O?�Ez�7� �\N�>�n��'7��dߝ>�С=��g���=z���<��[q���<�j�>-��?�|>��"�M�L>(�3�AW�<
��>�_%�^��>Zj�>4��=���=�?D�v?1N.>`SD�.2P=�X�� C����il�>��?��^�P"�=��>������8={x?=���{&?�!g���=���>vY�>M����p>�^G?�SA��=��)=K'?=� $>1�>�&G�Lֻ<�A���Ǖ����~���\	��x�>���=d@��ߋ>�5�<�.�7���B?��w����?�z�\��q-+?�Ӓ?U�n�y!���v;��?�m��k�v�� 뀾(E"�f:�k����0?�e�� �z�A>��|>��v>�Ec>x����ό>���>���Ԫ;>r�x=(��e(>�L���/��.>��?�վ�m��Ao�>���>j�����ݾ�����8��ū�JfͽSƾ���	� ?�s�>�mF����n�>v&�>,ֿ�ԥd=jX�>��p?���>�4�>/��Х�\�%�y�����A?�Z����>�!?ꇆ�rr�>�N��Ў�|t�=#�9�1���I��Y�>��>���>���=q����G�����R�[�S5k��>X�E?�&�>�?�M��o�>,x�=�ʾ{`%��>|��>�	>��'��?�眾�1�����1�?g6�>��/�B��~T����:�1�>ظ��] =�?�>�r�9,����4?�M�|;����@��ff����=�E[.���>��>&��?�� ?�H ��m��ʲ=�1P>�ݽ�H�9��N0>�>��d䱾��R>�d?��)>��>�~5>$�>gJ>���?\z�>l�ھ�ѽ��ｗA(�A�B=�y޽>����>Z�>k8�>��ѽɘN?�yY�ɖ�=���>,�?侽J�b�P��=�">YD�=6.���?��υ>���>�0��1C�����P��>�ݑ����>���>;�?u��>>��� �>�
=��K��Jd��6� sL�|#?p�_��/m����=��k<S<W?�B��-�<�>�nY?�C���WL>�?��>���>��>y�o>X徥F��eC> J�>۠M?��d�g�6�����Fu%���$�
n�>��]?v��=�����>ڴ�>��=+���+��=����OG�{ ��ë\�y�=�u*�1l+?�0޼���>#=?�ST���W��V�'�
?$>ЁŽ�rŽ��>l[l�euо�H��e'�>1(?�?��>~c�>�
����=RA?�?^xd�G�?A��>s��[@?�d>��>���?p��>Cϝ�� ��X>��<Q�/��q7���
�j��>��X��O�"?����L!�8���پ��9��е������I�TR>��Q?Qϛ>���=��Ը>-�`?�P�VK��"30�� 
���w�s�r�?��{>+eO>{78?���
�>
���ŝ=u?��K����>��?��꽏$�>�f*���=Ǎ�� �>���0��L1b=S����\��JK?�X���T?'N>�<���>��?Hnվ�,?��M?�O�=�V7��B�1���p���oJ�Zϙ>�YV��]�>3$ϽX�U?�&?�he=�Q<���Z�>\���V;>��W>�p_��j[>,D`=�M+��&�>)�)��qH���#<�����#��4�="����F�2N�>�M���Ք�A�1����h��h9�>l�E�%��p��>�;�q�=��->AJ��wl���2>w/>��ڼVt�=��]�a���6>�P?���M�	>�+}����>��k>��i>�Gj>-V�>k��>$落v��ZN�=��$>��>��c����Ũ>�>Ը>8�پT�I?��}? 	?����h��/�=��W�Zu�=�Z�4W����~>�NN��M��(>a�о@#$�Sĳ�nݾ�!�@|H>t����Z�*�t<O�>A�-�Ñ۾vż>Tz�=�g���?��C�d`�T>����c�E�4�|>�����;2�VCc>3]��'?x=M?S�)?O�>�C��6C>�%�>�w.��*��^��>fζ>d9ܾ�0�>��>�t?�>e�����$>?�x�?�F?�'��T>x�=���o��UH0�,R�����>���>�oѼ���=��>�Aq>��?&_?8�?�2ƾ�i�>hX��($=8�>f�?�jV>do{?��>Z\6���W��b>��[>���=�p�>���>WP������lt� �8?��E?=s��Zξ�%�>�Z��6������;?]V�>-��� N��=?��=�ؐ��1��x?�X�����q����>5侾�ą��=;ܷ�K㬾h�?�ɠD�G��>�@������
��.F�>�6-?&�;7X>n,�p�=�J��q�>��$�{g־�>���=����';��(9�> �>X����>H��>���>�z����"��å=*2��(?&p�=��>Vnv<�{>�������}8����=�������!��������#���2����r>i��>�1�>���X.?���>Mp�>��.?��9?��$>*�>��>Ҡn>�5�> �>��>>N?ę�>���>/s�=6B>�T�>�l�>�,n<\ɟ=ϑ��N=�P{=lX�TS��]�:�P�,�M.?r�N>`#�>ڙ�>�]$?>7�:���2��
�>�����㦾Qx��ގ�=d����E;�O��<K�}��9��z��4	�����/;�=mYL=>,�>�=�c;~���m<�(F��l7,�	¼���=` ?a_�> �>Z��>q5?�xj>���S�i���>j��������=�uy���@��Ӌ��Ƭ=J5$>X��>�&�>@߽�T(���B�>��>������[�B<4Q<���`b�����uJw�B���T6߾�S���
���C=�_o>`��c4>xe��?l��"m<���=j�C?h�;=�Ρ>%�l>K#�=�"[���ڽM�[>Ì�>�3u��l�=�+4�>�)?/y#��^̽�r��7�>��\�Z��<H69�e3澔8>����Ȕf�};��Fz�\%��G�>B\�~S=���⌾�Cݾ;zy�bT��"jL����D�BWQ�| ��	-�� �F�������F�>�ž4ɾ�]=�l>�r�;f�A>	>+=��i>���>~�T>m�I���۽�oz=���
ٖ>�\����=�ZP�Β�l����>C���?>��0>�x��\��XѤ����>QF�ӯ��h�ﾂ�>��c��ǽj�����>�rN�+=�>W����<�>��?΀�>�W>(��>�)=>���*�H�t�>�k�	���=�ھ��쾏槾tu�(�5���ƾ������>J��<iA�d�f������>��&=/ϱ=ĥx>�� ?g���	p>I�O<�fi=�y�<�r>��@?~�U���&=ʁ�>U���Yl>*�^ž�uܾ��>�	�9�8��k����>�>�N>�y
��ȾՆ=�g��e�?���9�>� >����{$�%��=�B<��>�����p�vń��1F�/me�JÔ��V�@?CJ��K������֠�I��˗���8�I>.;<>���>C�?�!"�+�>uO��e������=|��>S#�M��=sw�<����È<G?=]}��򨾉���.�=(�$?��Ἄ�1>QV�>ڹL��ǔ=�>H�->��R=HdE�����W����(���fk�>�]7? 3%�vO�=[Rf>%Ml>g$���q�bo>��=(p=�l���,���־�r�F|��a�`>&����R������$��y"�>�"��6��=�UH�:�=�T����>M�=�9�>D䁾$��t)��P�>\Խ�����a���`>��>�w>�`6>���>m��>o�>4e�>|�'>h��qu��w��#Y����M>������>PC?`��=p�=>7�>R%>A��>��/?�҅>�'�>��=���>�)�<��,=�V���?tSZ>��>h��8	 ?l|�>��Q��
�+��=��𽍕=@�^���_���Ͼ�S���y<�^w��{�>�sr?CN�>	�;>b̞>��P>�!�=�ť>��7>��=5�>�Z?Ȭ�>�����Q���]>�t�<��1>$L6�z����)�]�G��1��)�[��B�~�,�!��84�>�LX����>��ž�?���>H�Y>���͊>5��>Q":>-/����>�!=�\�=@�@�ܾ��3�Jف�`mQ>>S��L��x6�}X�>�j�R����@�R�>]���9�v>��4=l�>@$>���H2#�F��=M~>;mq=x(,�θ��l���A�P�����>�u���.��U�������ľbè�]wQ���-�ڽ��7>�V>����S�>�L�>4I>�l>��>��&>*�L���>ÑR>���>�m8�M��>'�����j�+Z���d��V��{��=}ѳ>ZlȾ��;��h<= ?�'�4��F�������ݾ#�>_�?�[�<�݌>e�k>�����T��? ?<	�>��p=��%���;�f����"6��9/�r�%��̃��*>''�>&�g�l�U>?�	>"%���Ģ�K��=� ">OPz��5;?��~>�p<]md?6O>ϭ�<�E�	4u�E����C�1S�����I��)��4*�� ~2�H?�Q���>�->��?�R�>��>$�����>J# >{I����=6^?�M�|WK=�|��!�R�)���LB�֓�>�T6���L��>Z�I>g���{��
�վt���y�>^<=�>x�ɾ��A>H���,���z�X��>Z
��i��=r�<(&=�׬�^0Q>D�?>(1T�f-�<�k>�0�>h�>�Z���>F��2��>�ҽ5~��wLо�%�>9�ǾT���o�ؾ��h>uJ��瞯=��=�4>e��>��>�c���tv����>���ڌ�����a:����=�!��|t���]T��&����5��>��>�>j�����k>�z	>��=^߾�&>�#�$�<OH���žO�s�gkľ���*d�ej?nt�px?G6��CO�>Jo>n2?\��8��>���>Ƶ=>��+��\�>	 �=��>O2�~T���0�)�>2پ*�V��B�>MV�k���,Q���ґ��ަ���=R�:��c�=x���>��Ͼ|��T'>�z>�@��-kݽź��s�>�Q���i=�?=:��>�P7>/)�>>�v���W=�����t�>�U>73���O�����->��=�U�l�$>�?��?>m|><�d=�"-?��?���>j��>��?�t8>P6����F׼��=��>�ק>;��w>��;�>!5>7{�=h��������k�3Ca>�큽�ʾߖ�� N�Za��Tƾ���s-���о��Ǿ��R���,���WD�>���EF>��>HТ>CW0�g�>2�=��=�Y��<���. �Ŵ�>���<��>��l�]-��!z�=���>9Y�>�G��f��: 5��:ݾ�7���Ծ�
W�����{�Ҍ7>�yF=H��>�u��[�>��>o��=������>�p�>>�P>_/���> 3=g��=,tѽ��>�?����"*���>���p�>sÊ�I"�>+>��"=T����a��賾k��\TT>�9z��T�<�EJ��"�>_7�P�;~���>�İ��n���7����<�H�*�=��̼T1��ݏ�y���:�4��T��Ξ=��?����E6�=G�j=�n��h>�w=lB1��琼�f��m>�˥>PLy<���;�jV>��5>�����&W>[f	?�_�>�ى�x	��]����= ���5(ֽ�\F=����/����豗>���{T�>1�F�Ш@>1��<hߙ=5؞��`>�����%>D�F>�������پ僷>4�����TuM�#	�>�^������sT��Na�J�㾐1�`��D�>�k� �@>K ����>gL��'vľBc��Y��>��������������K���#��M��j7�����h�'=ck?�����sgϼ�������ν��e�<�'Ƽ��u���ս�L�:\>�=[g��H���4~�ce�>Z1�������1u4?� ��Y�;�Q�=le>W�����y��2�=Cn ?��>U��>�W�=�
?qe�=l��ھ�!��-�%G,�0� >iu������#��W�����>]Y)><��>�Q��>�>�	>.���Rƾ��>���<�a���ޜ�Ռ�:
�ھKW������ET>�F�xZz�|R�ǿ6<q��A�	���>���c�zΈ��?���� >j�v�`�K��}Ǿ�����\z����B��,'>qO?��>Y�?�ۭT>�9<⍋<� �>��)>@ժ��	?��轄'>>�)���Y>R2�>��t�p��d�+��*>���d����E+�sŞ�Y����Խ�k>�*U�!��f>pj>�N���w���=2�>O�Z=���� ���>��޾�����"�������>�>��=q�>���=�^����>��=�/�c>4��B4>�7�>B>�X�<����1>�*>!B�=k�w�'��;�N����>3Ќ<����#�>:�>}:ϻ⍄�)�f��^ؠ�L�L>�X�=u���ݛ>�==��Q����h�=��j>��w�@M<��c�<�>��q�b_!=ܦ'��g��c��=��&>�f?[0��")�H|�q��>�wT��l��ǽ��>ꂂ=v�z;lN��6�>Ͷ�=�b�>_�|�t	B?7+����ν������>v9�=����I|��}> �>.�߾���<��=Z�>n^���a=Q��g�߽K�3>_�">Kek�{\����>6D>�ý���߼ ���Z�q���0!�>M���0�[Cӽ���>_7�:��I��%]>��q����2q��z��>`�>\H2>��s�H�4?h^T����]�=�M�>g^G���i��~��T>\~ڽ� �9.����>t�۽�˝>��<@�>��B�n�Y���m��!G=�g<����=��]�D�����>�F@>9U��"I�^H���s=�.��*�*?ט;KV���S�=J�>g] <�$ֽL9��h�>D>ZZ��%����>�V���:�=�I�Ô
��RB>���=tr� V�=%I�=ᆽ�q<ER��e7>�>�L �B���:�e�w�ym�C�X>*��F�[���>E�G<:24��aJ�S�'=A�W>��S��u��D�<�5�>x5�����=z�Q=$��=�� >	���"E�>��D�ϾY�t��.*>�ng>��Ƚg�0���=�"�>�-Ľ�]9=+���>��=�CW��>��5=oͽ��F���;>Ws=�e�*z�z@�=�?R��=]ʗ>J�y>	�>$����<S�=��<)�B�o>oT!�T�>��<�^�=b���۾jQG�2�_�;�����A��.�>Jٵ>K�l��rJ�&�>���=���>�Do�=��i>��><׆�Zzc>XXQ���;>v�t�n�C�^�=`�f>��w���M�Al�>3�Q����OYE���S>OɆ=� 3>��=�&>��!>��ڽl@���o̾6Nn>I=��7>���3�j>�>�a>҈�����	~�<�N�X����ɽ}��{���I�>X�Ծ�㸽YZ��?i�>�H��7�i�Z፾�q>3��>a�>�~><%>��=����b/����e��=E��=́�>o!��9���]>��>��*-ݽ�7��\Ϭ��TY�����Ⱥ>W1|>y���D��<��C>{�A>EQ��'��b5>w"F>�'W��4ƾ>]3��p�֙\�yU[>n2#=�����GQ>��=f�&���p��b�>�&��9���݂���@>B��>�ڗ>���>�]�>9�l�~;�j�G����k�>�)�>!V��������N��>jT�=�E=(
 �[0�=�t.=b�=�#F��Ժ>��>ا�����E>� >w� >^������$A>��;>����t,>w�� �h>�
���#=�U�<�}�Qj>E�}>0A���<d��=����:=��j>]��=�ɛ>(o�=��C>h���%>��{>�(?�Kܽ�T|�)��<�?�-�=*����{μ�@�>R�>fn?�V��<�՛��/��o�>�?�>���t�P��`J>�'�=��w=ߺ^�9|�<<��>�,�=/߬�yO>mY���=�\�>�v���W��2�\>�=y$�us0�΋={(?>�z)�Y���n4��ܾ>J�'�p�,>���<��=�杽���=�0�����>�m>��E>_ξE]>�b>��>k�hߢ��va���Q��X���h���ֽ�o>p���0� �!>��'>�I���!����<�]�>�¬�C�����>0�z�vV
�*��Bb��>�=��Q>��¾� �;�V��M�n>j��3ӽ�x��F"0>���<$�=��k>dwp>�#=��D˾O��T䴾!�J>�kl>tѼn�׾��>��6>��>��t���B�߸0>GL�=Ъ]�42�=�n�._=*7�[����ek>:>����7�l�@N�=*̔>[3���������>�<
J�:�>'b�3:m<�D>�Ύ�5�i��5>�]��l���ݭ�;8�ؼQX~�I�H:Q:�9g���	���/?�ݒ��Bݾ����>|�5�~�y��F���\>�>�>��W+���]�>E�*��iL>i�@�"�=���b�V=�
���4����"��b�=lLz�}��>��</�;\���� �����9(��W�ܾ~�R>��>'T�B��>����^�aP&�Mw�>`����1���݁���>���>6��U>	#�>h�L>���C�y�^L�>M�5���f�S]���;�Tu>p	��iN��0���Oۍ>�6��T�=�_M=pJ�=�@�=ҭ�>Λq=[�������A>�s�>g��Ҡ���<}�<���_�%i��a
��Ӈ >18�7)��z�Y����>>[>=Sr�:�y9�.>��=��q>����pCo�:�f��Ą�_-����'�嫽>��>���<Ia���p>Z��=�h>B­���˻��B>G��>�̾�`m=���k�g>�PK<�|W��@&����=:�Ͻ���)��=/^�z�>N%)>����˻��L�ܾb�&�t�����T=!�>&�C=���>�ۯ��p�<W�߽'v�=�[�=��V�{���[d>'+q>�rX�~f=J�>�6>�X�����N>�O��Q�������������>O\	��cb�\.^��n�>r�>5"=>��>�/c�!��>����eח>]��>�p���(�=���� �=��>�3�>7w����=�j�3��kP�=ܛ�>u�K��(��'EZ���=�h�N'>�X��W=�vL=��=����1���Ѿ�����i���p��r�>�k?�S�>�ƽ�C�:�I�^�.?h�#�l����<�u�>\�J=���*3��鵈>R��=fʽ=r�6<�1�	�=*�<�k6>Rd �����P>��6>l:?��2���̾����/:�7i���@�>[B�>s��s�-��r>��_>AL,=�{�� �<�>s��=�\���kZ> `����=�ϼ� �X�s>�2M���Ƚ�|"=�E�<��ý=��I���%>>�}��^o��Q|>	�i>�B��>�3������0>�D>�'�ټ��E,F���>��1�e������)�>�����/'<e�ݽ+�@��|���N>r�ξ���-o�=��F<ఌ� yI��^��a�>v�����p�>j��dIn�(k�E�E=uO�>��������g}�;��>�_��ӊ����=�3�>��p��᛾$��>H쐽��E�a����>gڶ>���t�M�M>�@i>�l!>L�� ?>�`q>t4O>�ӯ�����(F�~��<�~�>@ɾnmҾ�(>�>L(u�Z����ʽ��!>�6Y�4���Wh���>��o��:<r½9�>�Q����/>z�`>���L2�ʇ�=<Ǖ>@M%=h_m�,���Q�>綹�vL_��K������̀>�tO>X>]�t�0=��>���=������ >>s�|>y�>�m�
��>��>�������k�=��>g�Q�?�N���ýJ��>�O���h�Ph��*��>E
���!>S�M=��?O��>���.V�>���>[�����=��>�=�H�*=c�<cڙ���?D�C��=�ϼ��?��~=L��2�+<-W�>}���`J=�x��L��>T�]�O�S=�Hn�	C;Ϧ������/�3�#?��Ǿ\��i�
���A>�Ф��P�`�~� �[>�=�=�B�!XM�U�0>��=��u�<KT��Ǉ��_w�(�Q�|DT�mՌ>��>���K��f�>�0>8�4=5���W��>7>�|9>%����}��>���>�3>�E��e,�=�\>ԣ0> h�$q8��Ӽ�� >)xy��!�
���i��>d�T�m�y>Ĭ
��;3?4�$��˾t��x6���e?O7�=�B����#��?�i|���d�KG�=ri>r5�=j��=�|?d��>��>�;�!��?:��>r�0?�5�>��>�a$?@_>U�>K��>����4m>�͌?��V�D�վMC=��1>eU��W�J?��>�a>�=>��Ҿ>���t�s���/��W<�u�۹k?�ҫ�Xr��:Ǿ��=ߐ�>���
	��Ҿ�z$?�d��W޷��߿>��--�=ʯ7��?_-O��K�=׫ >�L4?�	f��_?
��>p�̽;�1�@�쾶�
���?���>ޭJ>"���xc�?��(�cM��~��*?�Y>#�j�������>gx�>^@I�4(��l>rBb����Oh�>���o����\���>� *���E=٦2?��>AIB>y@�����=0
��M)���>�l;�����W�ڶG?d��=6���8���΅��)>TlS��{B��Ȁ��w5?�">�ߔ=�N�>����Cw���>0��>7c6>C�ʾ���+�>6��(O�����Ì=78c?[O�3�T>����JӾ�x>,� �l�=�>�Z<�<�^X�ܴپ��>mw�>ݾ־Z������O��Q(�����>�e ���[�A�k����>��I��#��rݾ`%>2I=�~b����ྱ?�>sӢ��k@=�!=��;��|<Vv�>@1�	����7J�E�S>\��>�Ll�ǰ�>b�q=��^>M1�����C���h��H���3�tt���M?�mD�<Gv��=��n�>���>	w��H'������%'?� �$���8	�>�c�=�=�e�>Z�'?p齭���+��52��A��I�y��	�|�>�8�>�<e�9�>�~�>w�Ἣ�G����}.�>�;�e޼�JU�\W[=��H<��߾�Q��gF	�A�E?��<Hv7>��	?��_>j�=#t�>܂ ��<�����:�J�Mq��~�D>���>�C>8���K	��Q8���F<ᖢ=4ӟ��|x=
T?�h�������V1�S� ?��<n��>��>�U?8C����۾�����$��tN滖�Լ��[��j�5��F��>#N=�㘽'�
?�y�=*6���ϾH�*�Ypؼm��>Ҩ/=��D=.9?&9�k�?ij�����>Pqk���f=�>F#c�X�o��׿����>S�_>�������U�>zL%�\�?M&��V>϶�j�?	�>�\8��Ej�#}�>t��<�y�>�<=
�^?[��=�N6=�ʅ>� �+\�=y�`��j+?�o�S�j=٪v=���>��L�*7���=�>�)�'l"��?�>��>���<�K�?��<���<�~$?����	�l�>���>���,}�hu�;�$=Z���c>�{�� �	�\L�>G\νu��x�<`�>��!ؾOoM�ˌ=@�N?���>�==ܗ�>��=��kXؾΞ����?_0?%L3>��!?��&$?���>��>����wX>���?�ʾ�%���	>�JF?;�f�)�/>a~2=hA?��>�i]��^>TM=`�>��y�>�@>�3�>���V�>���>]"��Q�?W�>vƿ�?.d$>�.>b:�>��s?_�N>p};��Ŀ�,-���Q>h>M�?Dpa>��Q��>��zW�¼�>|`��T�5?M��s������߽��H�~����ԇ�f�>
7?N��
=���>�*�?��>86þ�y|>���<_>KV���>�'>:o�>[I��$��sZ/��<�>�ͼ�h+Ծ�ƀ���Ef> �c�r>�F�D%O?z�2��/����<�@�������5>Z^�f�<��i��K>w2o�a�?m�+?��>�������0� >밾��z���#�����k�<�.����(>jWH>�D�>��1��;�>�L��~�󵙾�R�>?��>��������
��>��;�w>�����=�	�D�h>NZ��/�f��Ɨ�$Sb>���=6���Sߚ>m��>C�b��Cؾ�f�}i�a��>���
i�>R�6�hh?'^k>U�>1p޽8�L<�s:��ؽ�*K�$��=�4�ؐ�=��uu�>��n>?�w>��>X��@�>���=����駾AA�K&J>�㍾<�?1�W>�j���B?I�/�M'¾�&�=�8���>;r$�PH>��=d���f>j*>�����X?�����_���}��>�Ǜ=�Ǿk���ށ>m���e�=���l �>�W>=T[>���)[2�l6���x�;i�F�B��n���+�oV�<�"�?�&?�-}��R��O�H�E����ܺ�Mr��9y>L(�>:t�=<R7?g�t=�^� �N�w.?��_�����ʲX���>"?��iT�4�9>E����E��w���&)?Q��ۣ���&&�nA��S��>����8�dC��0�]?/�'�/��[�>/I[��UM>Go�?�]�>��A��V��̋V=�m��m���Q�G�LH��~g>ۧ$�R8�Xi(�mâ��;>��s�2P�>��߾I�L��W8=�����쟾�w����Q?�L�>��N���񔽫+��\���'ƾ���>�/V?�Z>44�C�Q=f�?�9?�5�B�=��<6�>c-���Ev>�=�?�r���۵�;��d󀾏W�Z������>��e>O���<>:�>D9�������F����=�.�>��&q>����^(A?�0��l�V��
"�mb%?��ӽs�+�H����>?=վ���>�?���>\�=lFݾ���>��?Y>噉;i�>�C*=�Pt��N���21�[K>T��>Շ?��j?\��>e��=���8�o?�T�>+�>%m��ϻ�>�>�1��#��v��>4��>�?+az>�1��zd>���������4��ωɾN��=Bu���w>��??�P?K�����h��s�>l$��
+������/�>(�H>�?s,��%HQ��bC?Q2Y?��뾓)G=&j�<���>D}��2A���R���%?Lp >�!��?��Z>j뚾��=a��>5��LO3?�:=?��>��}<ҍ��t�=h�����l�W��=�w#>��#?�������<��?]1�?y�S><ܾ���=Bn�=\YH>w�+�;P�>'��>a��>ɾ���6��� ?z�0�|aF>�L>��?��v�x����>�1M>[������,?��Q��I��M���k�E����[�>D5��%�Ⱦ ����"	���>�pB��ɣ�������d?�^��(��;C�B�LN�B_#>ua���W:>:0+��8�>����`].��q�>y3�>���g�� &�՟W>��N����<?"� x?�f��4�>��b>��?N�龻R8��@?�!������G�P��1�>�^�>#���҉�m{�>�H�>��>�
���ݽ�k?��#?�N>��G��>�?�x�L?־F��8W=Z�������~E��J1>T2���������������c�>R�,�K��<K�%?*2Ҿ��m�d���]:>72�:�#U��w>BMY������j�;����?_����d���ȾK ?V�Ѿ��	��n���+���H�����T\?��;���7mо�ږ?$f>4����[���7?��>c���J�?ؽ*>�\Ͼ9Pa�I�i>�w�=�hѽ8�徫v׼X�z=�,�65P=��սV��>G0��5.�=�׏��;?Uu�>�4��N`2?��>"�Q>L��.��8�=?���m@�;�>	?e
�=���=����G�M?�  ='�G��>kr�>f�>�jr���a7�>����� ��U?�
��>���<�↽��о���>�%��C�[�%3*�ᰥ=x �=���L�1E�>��=������Ծ[�?�[��Q������E"W��@��p�ʾ$���g ?;Պ=�B齿�J;JHs>:��>�t ?��Q���?�5K��@��|L=�n8>[S��.�}<m7T>��Ѿ[&�>F����!?R�s����<����>)�0����<4�n���a>��ھ���=Rc|��Ɖ��Zҽ��W=�˾A?�/2?v�X���]��������>v��> k�#�W�ﺾ�^�?{-�?A��?�𳾣��>��>���?71�=R,>��->�*���>�U?�*>�\>ɾ�%�>�e>/-�?���?�M����>�k��`�?l�a�	�?%K`�!�.�R���������ķr���L?�뚽��{>�f�>�0q>���<�>P�?�����x�>���?������<�Ʉ�����k翲�^?�-e���a��*�?[P�=��>����#���s��?���>c�=�3���T�?�턾��?Ru�_�*?%��=7�?��|>���>�4?
E�墾�Cp�)X$���h?�Jz�(R�=�g��Y�����?�I��\���6?�g�?��ξEظ=?��>h%���r���(���N�+A�P�{��?�<;�}c��Nؿ;r>��>�:�6&��/�پ���>ɻ����?e?���?6L�^��	���u�z��I^>!�qN�>n�</��Y
?��?�w�==�����>�M��b�?���??+$��ڟ�<u�����?6}!���L<�ܡ�>�����>����9|�4�-�4���q,�Ì �<�=��׾����_>�?�|�������$���(=�����P��_���@A?�-�>��B�R�2�j}���ܞ?qS?��H��x=o�2?dL?=i!�xߕ��^<?�{��j�B?hW�1$D�R\Ͽ��+�����C?^�z�x|?�Z�>~����b4��3>?@h?%���{�L���e>���=ꋣ��a�����MI? ��=�V_�x>q?o3(?Z�������~��/�?���>����N=خ��ǆ=��r��+�>b6�> ?�	��;�v?��>%�������[r?!OI?��U�3؁���7?=�@?�@ý�]j?q ?�':�Ҫ?���}C?��������=�=��?(�ܾF]���'���Q���V?^弾��h?G䈿���JoX?�>:僽�Bo�9J�?���L�{�,<S�͡h?�\>@�	?����	B?Pb��B�>&G�OIY�mW��Uݿ���>[��=9�J�.F�>u&��~�>7�i�AF�>{�7?z���������>��0?��l��/�?�M��y#=U�n���?p6���~C?6�>E���?q>�*�>4�?��j��`�?d��XzҾ��>W�ÿ�J*?��.����������aB=
�c>T�b?}7��Y.���b?�U�>=
B��V��x?����>a�>aT���?𐿏N�=�Q�7��?\o-����q�n?�v?uO�>62f>t%��W?!�v��pd>m�*�E<�?7b��vr4�2��>�N(�����$��V��#=�+��ѭ@?�^�� �����>�ǰ=�.��Ӿ���?B�>�h��Ă��L��-Hc>�e0?�~J?�u>a5N>�F��>;?2�Qӄ�|�5?��?Z��>�{߾c�?%�=�9�?^������ܻ?�oq=�V�>��P?�?@=B�S�>F.^?K�?��B��+��?,�>`�C?j�ݿ�)̾LY�>�ʟ>�}j>��?ʀH��P?G
�C��=�)�>�Օ��9>fPJ��ȩ?/c0?M�>�L�3QĽ89=s.���m��o�r?ySU�ʠ��?Q�H�VT�Mr�~}�?"�>$jr?d��>�T,=PD0��;Rru�+� ?�ڗ?�󮾾�����A?�$;??�V=�>���>�{>�g?!2��1�?�Ɛ?���?@)?�;E��eꩿ��ɽ Q>�S��y]2�?��>h8��p��,��pE?-Q?��.��Ծ�Ty�Z��=r�Z�z��=��@������=�H��^0]?��*?ʈ?\�I>�N~�4^���φ�^M����=�¿�(>ݠ��!Z��d`	���?���d�X�?leF?t7J���b�����A�P?t8��E�>R�L?^�O��V?�q>� �ʚ�����>�&���X��c����?^p������s�O@�?�A����[*�dCx��o��xG�C�5?�r��0�;I�־A�>�ū���>7�?�y$?���/��?�JY��bټzD��0%�u�A��>�G�����L�?V�i>����ѩ=q�'�	������i��?�t���=�ܔ�M�̿s�F?���>�㬾��/?�M?(���>; �s�Ͼ�T>s�;w��?�@r��*��)��>�)l?f!��� ������?�����|�^?�FS�{�[?''�U�`��v��)t�;�0Ͽ�7����>��+��?���Ì���2>#$b�$�>x�/�Z*�=	Q�<��`�3,-?�1?�Z�=�w�?�����=��4�� @��ݽ���39�����>)�>���=���M>jža�q?�|��c?�3�>��z���C���?��?�8���O�&U?ۄl?���=��ƾ��z�֞�=�??U��b��?� ?�o�>2彾�=b����Q�$="6[?w2�=��>$����M6�����j�%j�����?�Ԯ������N?�8��P���f����?:D��^z�?���\(�7��;�%�ccȿ�,�?a`;?9ד�A�����?�R�>ߤ�a 4���U?�S>�+�>`�>���?��?�B�?��,f�>�������17��!�>U��?C�a>�W��wᾨ;�?�'�>*��2>�>L1B�-0?qa����?�b�=�>Ҿ֒
��l�?�;�< ���GͰ�}1Q?堿>����󾊖�>�:k<�k	?Г��JU=���ƾiV8>lѿ��f�?��!?a���ě���
?�ك?Za#?���=�>��)?X߭��Z�?r�]?n9Ľ��!<��p?@/����=+=\	�>��Ԛ�����?�}���Y�=��3��;h��	5?����>��ky>��>AU(��
=�P�7?f;�����	F��j�UG���7��p���?d�?;��I,���\?;j=�Ď>�Z�<�*?�+���W?�F�.��Ք�U�@��ǿ���hX�>��?�F�����?��?��	��Z
>c�;?��?��l��P?�]�y\F?�朾e߹=��>On?�Kr��~�C��>+6>?��ٽQ>��)�>�@�:A?�¤�\T?9)�?�? ����뼾Ǹ�?jQ���@&����?��?/[t�ih���!>#B>�M0>z#>"�?�ֻq����a\�"�;��n���"��&V>(S��+=a���=����WI��9����,���?NJ���3�ECs�hr��ʬl�O����徾7�>;|.��!��J[<��t��f?:$?�].�Ҧ�>��O�CI>����x����=�.�>�`�<�>B���?C����#>��R>Ԣ?�����;����?D�I?<����?n���sB?�{��L.c��;>��=����]��S�>"���-�]?H=��Y?H`��z�uЭ�{�ž�r���S>U�=w��	B�x����P־�� ���c=�ӾR�D>)�,�U��?�����`����������R?R��=��S��6�>�����	���>���>���?
�����X��>���09��H���P?�"��&�>�f�)G���\�R�&�/���赺>�:�>(��>Քf��m�>8�?uN�������>+h_�&y�C<f�N��=מ�>!�>�ˁ��Z`>2t ��y��Z�=�媽��*?u0>����j�?�n�?�$�=-J2?Рƾ}�X?V>8==�?MG�omj��
7����e0ɾB��>~,�>:��i�?ZZ?H7��9�1���>b�?^q�����<�񶾊5��z���F�J�	D��Y���1ȽhE��kg[��G��+=�K�����,�,ӟ�}ɭ���>>�O�v��kh��n
�=��οW�D>e}���S��z����6=g�L����>���>���>��پ/l>�2N?�Ӊ?`�Q����[ 8?|������=�n>�ӂ�b�.��6�>�.>�v����=}���&��G�XR\�J�x>Mw��	�#?���>;�>��>��=���>7Ym�2:��|.���5?G�ܾ!�����=~j>7Ͼ�,�X3���>x�G?�g>�e�>��>��~`�>'32=�iY>�B�>�MR?"?�f?�d�>�k���~�?p��<��
?��d?��H?Tl$�bn��3Z=��_��zH�d�>囍>�Q"��y��[s�)�)�wq��24>с�={�4?�>?�X�=��ž���������>U���*s<��ծ>=di�_	���$s��<�^>�N>�͍?���?Z:Ҿ�c<��D���?]6=�{>;Kѽ��>4襾,Se��ϝ�M��>��>�w�>�S@?�s<?BC={lо�(���=\�>'5;�J�1�Rn?n>�<"f>j�d�3>��a��BN>���>0�>��Q��=�����м��>�t�>�p�>�����޾!K��>nk�n+�����kG�����%��>񥸾�qe�t���h��>D�p>������<Js#?��#<��U>�d�>�H`>����<꾸,��@^f?�c�=�[S�@�8�=�!?����+�S��W����7?��ܼ��>��ǽȈ� �Y�&=�J�%��ݣ�>�:�=3�����1�>��=*��A���~4��S�>���Rʽ
���q0��侺^>��R�F���H꡿�{�=o#�r@�����=ξ?�
6�s���i>�Z>̎�=��:?lR>�qT��¾q�]���+>�h�kL?a$�>y�*g����Ҿxf����J�s�>XY�=X+�>�k?� =�zľ{��
ة�<��>�$F�k\%�`��>��L=�JܽV�_���>�D�>��=���>p��>Ͼ?��=bz�֥�<��ཱུO��w�'H�>_f�=e&r>/�>���)�=��aޛ��
�n�$=�I��p3��ʶ=�u>�ƾ��7�	��>�U�>䐭>#�g�cn?�|н�R?踲>����־-��=���t��)��>N&�<C?�c[����cAܽ+n�='0����b�/��>|Q�>�y�?�뵾����=g�>�NU��8?�AY?L?�<Ղ���">ڴȾ0�g>�>#J���<�~T�>�[�@��.�&��E?��v��?�=� ?���PKE�ӊ��l\.�s�>z{�;�|�=�-x�Ɯ��V�=lxr?I?����⾯����p<��N?�4���=��#���>&� �fa��fw��SJ�=���=�m�=�ʾ���>(E>����C��=���0�$?��L�,��>&@�2�9>�������.	�߫����[>�?=�>Q)뾙
W�]n{>��q?A�<>_J�=���rb�>�;��u�>�Aw>����'���c[��e�<�۫=æ�>����/�>�M?[�[�x닾����f>�{Ѿ�V=byY�����y��\�=���[���9Å>�v�ǡ>�
��M�>4� ?�!?���`?�������g�f�Y���'������J�<�k��L�o�{F>�B?Y�=�F�>�ߤ=Q�νL|�?x������>�>�2?�N����P=���>6��?������T>>k�>����4�J� =��<+c�=����#⿾�"�Z��G��TF>-K�=�> ]B>Z}=�w]?���<��t>�E�>Ѕ#��l?���>�?�n?\bb?��M�eĵ=�J�#��>�����Ӕ>�z�>��;9"=<i��"Y��	B>��[�9�h>bY�;�\ ��!�,��=��>?im4?븖��ƿ>�É=r���O�ξY���
��>�.���\�=��Y�<S��>�]U>S춽tP'�e/��y�O>,ྺ����:�>�a�>n�����ٚ>�V�>�h?SA�=����X����=�L�>������>��>4�?X��~���IQ����>�9=���F��4�Z���0z5�v�<A�>a�>�2����V�=U�?�K־@X�<��=�'�>W�#�EA���;M��o�>�V!>8�@>_^|�G?�kO?�\Ⱦm�6�^���6?��j�>XB ���U>U �_*;���9*����e�>ɩL��S̾^�>�R?Xh{?7����>`A���=?��8��O�M}�QqT���7�68h=c�1?2ߤ>zO�=�~�����>Ҙ0?n�"�(岽B>�Ë�>�z�9i�>�J����7>򻋽m��>�  >�5�>��߽�V9�t|���Ry�(H~�X�<u���>��	����=� ��w���X=��7\�>��>>��~��.O?�:����G�{�Ž���>G�G� �>���g�>��> LV>�Fʾ,ʁ�����^��d�J�ӞV>x>݄>:i��+��z�ԅ":u����>)e�=���>k��>�?J>j���Խ��(?�Ҿb�:��S�K��>|pW�&~�>8�t�^S�?�i�=�t�>�J
?[~ ?,]��f���W��b�@�>jm�%�Ͼ���>�֥=����<~��>�1>���>b��?��1?{�j���> N�n_k>����	*=���=Zs�����x���1��YֿK3�>��h?;��>("�=��=��(>y'�M��y�>�c->�?�7,���/<���7��;H�����#��;ݖ>u� ?
�����0?�$�?����+��>��=f4=��C�>(�<���3>P(T��[�>%�?�x>���J���B��N;2=�c>f�#>+�>�� �X�Ҿ��
�>���;�>������=�@>�!�Ⱦ����?\
����Ӿ$���ۅw>2(�;��'>p��nU�?5u?>_A�>GY��c��	8>t'��z��I��>Ym�>r�D��d�:�u>�MO>U��>�$�<�3?ß�>�����=��>w�Z?���=X&?h�&<U�e��� >�'���	?3��>Y�>X�=�,�<�ӿ>*��=�n�>��;C�� �	=�;�]6��utH=Fʁ>�"�Jy��!��<�H��BQ>2�F�B\>� s>a�s?}�?{H���I(��m���?`>���<�>eڟ����>�Ü��l1�Tz���5?{"0�)&?�+?��$?쏽���<� w>��о+?w|F?|r>�nS��Ԑ����U�>�/�� 垾�̠=��?���e�<"����W�B?�L
?肰����>�ӯ��1����ž>��=���><H��mc��^���@�S1�� 8O���(?�z�<�5�=���;�=�Y�?8�AW��d<>o/@���T>/Q�� Xa>�`�>Y�?"��=��!�)����>�����Ӽ�J�>���>l�(�����ؼ𫅾$ģ<�|�d�Ͼ�O3��&�>�� ����=��/���_>�eO?�?�h�8�[��1s�>)�> P/�U�=�5����V>2�#?�Y�>.U+�u]ʽ{;4=��5?ô3��7>$8W>�5�>�5��Q����>�F�>1�?7x}��7漤T�>���>Rv�d��>�1�>��5>N�%�t5,��=��t��E�=>��R��?`=�'S>D}�>ؿQ<_J�.�4�_/6>��׾�3�=x��>�"�>��'#۾�&�=�L�>�/��2�>:�2>"7?�c��#�)�.���>1
�ij��
�>�>[7K�l3O��'ƽ�tN��)b>*��=��><C=3�E���w>�� ?�j@='�<dJ��b!?->��kw�>�����?V��>�`�������=���>�Ր��ܧ���[��>�0ܾX��$]>�h+?}�T=呁��q>Y�?�j�>��>,o4? �e?�9�>Q�>K]����>�ܜ��[����>vW�>��&��1ὑ' ��]?$  ?N��>r"[=���>�0a=Sy�u����$i?�(��x�=hO����>�����>�6�Ĕ�=����<�M�-⨾4J�>,�=�� �X��N�R?6��E�ȕ�^C�>��E�!>µv�����8��Hwt��֟�ۻ��ε>
ኾ:��Za=FNC=�A2?\��Z>;�Ľ
>��1?G�c>�L?���>)n�>{��>���_n�>���<N<T�ٞ�=�G�q��>����>>��7��=�$�Ӈ^�o�>�g�EYþ�'.=]�����!�~-R>�h����D�>g`��3���Z?]�h>�5Ƚlz���k>ì�>��?�1t=C7W?�k>��v? �M?�o�>���>	{$?S���N��h�>r��=rĽ�e?���6�>1��=���=W�F?�t�?_!m??�?H��>�վ����z������V(=\y�M$!?�g>���_�C�"�x��=�?Q 2�ç��k�=�/�����>J�?m��>���<Z�̾h�B>,�?Nِ>��繾��W?��}ԾS�t�׺�>�Fw>D��\�?���?Oz�>0CO��=?���>r���L�9m��V�?e�??�)�`YR>0�t? tľ�,U����Bj?�����>�=�&�>�#>$	T�W�
?+���@?V>��'�o��>C�>��оD��0�>Q�þΌ?$����F=������#?b�=��a�~N��.f�=��/�fڑ�0|�MB�?����A�?K��=�K��X�p���
�W�,�>U�}���ľ�dп�]j?��V>�WH�#�����>o�׾\>V-�>�6ھ�d8>�b:���z=�9���
t>M�!����>�:�+I�>��S=j���-�;�?�����'D��y>�J���U�>�
��i >Q��=�+��� �
���<�O������>�?�t������e2���M���>�ߵ>]F2���=k�>�NN?��Ͻ��"?��>���Q��8���ts��^n��0	J��C2>d�u?�+}����E!@�����(#�8J���w�b�(=��H6�>&�>�d>���=�?O��>�O>1���� �(a����$�q^=�9�����*?�e��8q ?�C ?��R>��2�;lռ��ľ���?�ϯ�R�;���=�t�����9���8��.i�>�k>'>'�>m@.?�ʀ��5��-�?ԫ�>AI>{���k>֠�����>�Ұ;?��>#���C��>�t�=_N�Tc&��k[�;�������ҵ=ͪ�?査?�Dܾ q�>؏*>�Z�>�J�]61�<��>��>?-���GU��|.<4IB?�EX>ͺ���a ��!�>���MY$��$�Rc�����ީ>9zt�P��?	'�=�Ą?>%?���@�>�rM?��ɾ�j�=x[>���>k�?��*��f?�*�>�߾��U��6?�����(�>�?S�E?a2�( ��Q���?���-�OM]>��w?g��>�c.?�_�>E�w?�P�>q�5=]����p�>%K�>Z�y���?8Z}>�9�>4&�>���>�끾5�>��c����͌>�ڒ>h�>����d�l��>D ?� ?,v�>Q-@?��N?EH���l=��$�@���]����B��rI�&ƙ<l'>�"�DҜ�8�E��D-���k=|/��d�Q��ܪ�>XKb?�@���?H�}�31?Z��S?8DQ>��H>�Ԃ?$	@>T<�>�IK�q�s>�aԾ)��?�] �1�>P̴>#t�>�f?� ���?`ꗽ;}��A���b?��>�
&=9�˽9S�>���>�	�׆>k�-?�/F�����4�>�kR���o?zYb�53h?�r���>>�����>����\�c�̾+��>���?���`l^���V�:c�?�r�?&'��)t�����17L>ҵ>�:���侻y ?�ђ>9��>��(?�+?�U?���>`�?`�>>�1ݽp�!?��?�ӻ>X4=е��'d?���%>�7?��?�N��"+龰�3>��=���|�}�۾��\�s����e����	U��/�Ӿ�� �����K��G^ؾ+b���Z��r��D����7��?��}?�rؾ�/�����Є<��\����=Ɏ�%��=�%��7�JC���?H�4��cb�>���?��?��L=J���%u��~?J�u��?�Gx��j������ ?U˝�y >P�?>���ih���/k��w^?��b��վ�z�W��?���o�>)菉��s?)b���־� �>@}��bjG?�?��>����PG��C�>��>~��]�@XU��dM��VJ>�ٵ���r�z�����k��Du>�dB?j'�>T�	�������>�B�>1|�B*?L���|>"X0�Fa�k�4�4���&fڿ�p��yß����=��W==`?�d>:"��uՁ��T(�{eo�z�>����?�7׾	 �Ry��V��y?�e��/��B��>���V�����=>���=/ >�>�r��K��$%<0�����>���c�>*�>'���(���W&���h�9����>:�$�ڞ�=y��>Jo�9��5�㼴m?�V��`�������y��uE���q�>�����'�%g�b��>¼>�a�j��>�3?��(�����6��u�����>�`��e;0�pJ�>��@�!U�=�K>�7>W�>����l�tڗ=&�>F�%���^��?�;~?"��=DA>�V=�W'����=`!{�ꍅ���H�(]�>�ip������u>*��>�j�>��m�uu?_�<�#?��z��=P�p���Rؾ{��//���=�.$?���?a�S>@M�K��>�ua?2���Qr�9>��>�����<�?-��>��l��=��>��?qq�>���,�>5��>ul��V�ɾ����V��>w��<���=�O?�/F?�h[�D�)�=H�o���W��:o���W�bA
������;uH�����?d~,��8��� C�]� >;>�q�>˨��]�>��F�0��\�"l�<-��Tpp<�U���h>뷅=�?A܆?ҫH?���>0�>��>���ep�=8q��7Lb�l<�ID�?�/�?@1?�?�E?F��>��<Hܛ�ƦB���}�շE��8O>�ů�;1G?r��>E$	�ig?L螿4�>O�|�}���h�|���׹���L?�E�>Z,?���?��>���#~>��7?f7R?�J�<��I>k�z>��f�5]Ҿ@��?�G3?�x?~�H��#������7?
�>�N���D�?hL�?�W?=���? �=i���&��>? �����p?�>$?#�V?걮��g�+�?���?]|�>$4M>��=��B?҈?��J;>�HQ?F��?]9�>l6?#�ξ0 Z?��>�u�>'�>�9?,�=҆>��W��������>��#?�1>�r�=�C���3�)�ſVM,>��>_�@������t�����0��A���G�RW�'$O��۾��ž(��@���'�?�>��<��?��ν��A�+x�j)�>�[ ��U>���,�Ⱦ!5a=(�Q?ڼ�>�i8?���>ŀ�?J��>N??�Z>>Ժ�>Z(�>5��>:�<��G�>Z�D=�ws?.z�j��=7��=`��>��N?�y/�W�><��=�Ѐ?^~����>օV=�yP?�}�q����+>X4?�Cr>�O����	~����>�y6>���:���A������q"W�yo���]?w����Y�����$�>�W(��A�� J��ž�j�=M�m�����I���Q��ۼ�+?�E��uz>�^��z�e��=>�d��Z�s�F��=�5�:���]���{F|?'���3����^��"��?��y�\�J�A�a?梇�T��=2�����|���F�fV	�+ ��𻰿`�����s>�
����#>�IǾ�-?>���ی�<��>�M��Q��HJ����>�[�>��	?1�?}��>d�?��4?�.�>��=m��ܸ���??��?��>��>�~�ա�>�p��ϑ�<`m=9M=w��?���巾\�>D����
���^һ�W}��p�=6P`�M���9h4�����Q�Z�D[¾~FD�e}?��N/�FV)�ԫB>�Pɾ�"�̴�����>5����+T!?ʦ�>[ށ>�t��xݠ<��t�)�?���3D���6��ς�����?n�Z?��>�>�>�y">z���|����b}>T�?G�н��ľ�����?�r�ڔC��׼<����$�=�<z�0�5���=� �=�c:=?&"��T��/Ʋ>���s�;b����>A:��|K������I�u��=@��W�>=�\=�Ⓗݾ>��~>R�Ͻ�C>�:�>0��T�k>� �=~�<({¾EO���^���`>��*=D��<�C�=&sv>U��7��=P�>>�X>��=#�G�a��N����r�0�=|��=��0����>[�:���>F7>"FX��aP>��(����̻*���\>�m˼���1D�;i1�a�<������>��h���Ծjǁ=�L?�S�=?�<�k>���>R4l������=���=��9�3^=�K=��}?}0��0��]>!��
U�<5$���=��-��!>j���D;g��<>�>F}��n.�>@g��NR=�#>���=p���F�<OW�>V��>��I>S���G��0�B��:W����>:E��&�{�۽qk�>L�罪�����˾��v>ǀ�<h:��;����>��H>le<#�o�N��>�z�3<%�f�k��>���2�q�)����o�>
 �CǍ��C��i��>�i>���k�j=�'x>p���pm>��
��è=���<�qػ����=%��=�e���>�$^�om���n�j��=�>Ṍ���W�����>�R>�3���)ھX�J>z@��,����վ�ǣ>�&2��&��Ćr����8�;[99��������DW!�s��=��/>�t��P�>�1�>߃>����o�3��H���V����>�����=L��m�>*��}��=,)���V���"%>?�C��2�����	,n>���\������=�(�=�'�b)*>#�U?�p�=:œ��;9>+��4ٞ>�����@��!Y=?�v>�&����B���>��>�U>�䳽�><�m^=89��{����>��ܽyu���Z�f�>�
�=�>+�#>����vt���c=����J�4>�<l��c-���\�2��>��H=rS=��	>�`�� ���{a���
��7���a_>�j��B���Q���2��e>��?5�[��`�=-�>�(�>H�{�8�>��;X�}=�⾽e�U��XE<k?̽Ձ=���<9�&���?O"�g1���rG>��>�(�<��	>���=��y=�L��l�B>��Ծ�Q�>�t�=��l=���o><s�>���B�W��oǽ�ϲ�#����E��*	�<4#�|�ƽ���>�΂�l���PҼ��>Q7g��I��&V�J"%>�>��>K�>z�>�=�T��>�����݂�m�j�m5?>�b��V���*T��vL=�!*=� S�$=�;�=*��=��c�S��{��=�*������	����<�;��$�W�<cS>�
�=�˩�����:��6�Y��8r>gM�:�����o�>YU۽M�ǼF'��w�=>'�9���𗤾��սb3�>5H�>��>�Qq>?m������)�NG�x��(>g}�=�-!>>��� �,>$T�>��8�n2o�a�=�r�=#�*��Ƚ�a-g>�@�>h�o�LtO�n�wȕ>T��>_r��N����s@>7�>�����	>��i>Ę�>�н1�X>a�ͽ����X>�|��>6y��&?m��y�<��=}Jr�"t>�y>�}>��>i`�W��|�0>G��=p=�����=��>�%?=r��=�
/>(�!>�7ƽK�a��R�<����]����+>fe�>0饽|�0�W�9�am?>�$>B�U�ߚ�=&�=�}(>�ɏ���=�B�<˨s=��>�6�C����$>�C>��>ܘz���{���D>�����<��]�8ݕ>Z2����v=o&=BK=�y>���=�򌾷�>��%>��n=a.���>��>B��=!{׽�"W��d<��J׾�g��}�I����.j�=��-�~=S]��!����=����:�=M���*+==}�߁>ׇ�=�a�.�=�Ԫ����=��=>z���s���]��]V�>!��������"�Ȑ�<��d<D�=��>HF�>SȽ�����0K�����rmj>�>�&Y�M�%�*>k�n=i�H�~ս���=�+�=C]��<�>܃)�L�d={+b�30�=7�=H+�}�<i�ҽ��f�t̠� 2�=��7��C@=�<>_:�=s�<�[��Hp>'9�=�@�A�?�F
�=�h�P��>�Es=$ႽYf:=�,�*f��T��-�= ��>p(�'">��Y�}f>z�>��9��M�BU�>��F���\�,�N�5�L>�Ƚ�b��0�����r����6=���X�=��h���4K<��>w{4>|�<�u4>��ؾ���
�!���x�>>�J}>���>�J��}��4��yY>�8��9f��D:'=�K��n!�>T �#{�>�8>��!>Ƞ��8��+��>}[�<��$>bR��Q��>��L��}�=�+���D>?����-��.J>R����>@8v>��H��I�%޼=��/=�l�� J&�b���
�>�G��ܘ�kr�-,A>U�1>��Z>��>��M�X�M>n��=�R¾�9�w�>�U`>0�Q=��W}S������W��R��Hګ��>XQ�)&>=捾�`��S�>6M�>�k;�a�=��t>ޑ�>L�۾�f�<�{�=��=�D�R�8�3`B=r?��o�=Fŉ=Ѷ�������Y6>��%>��C>4�>䩚��j��+��ݽ\�Ƽ��>���¢�>]�Y�Bs	<坊��K
=�5��߄�������/���U>8���q�>���=��=�n=:��ԅݼ�'���U���=x3�d��=6�N�ᚾ�y(�&�>"->�ic>MK8>|z=�ʐ=�󗽙�C?�#<H�U����>�f��RA>B
�=�	�=��(�� ��8�,�F7����ƽ�-�=�f=�ޮ=��E���%�{�k=�����K��G�>ץ�=��0�%V%>��(�α��X:���;�i��.b<<�2>腫>�T�Q���M>��4?�w4�.�=J�>;i�>W�����4�3�н1�m=���=;m��Ժ=Q�2=��=��=/��>881��>�x>1r>�#>J&l�O��W,8�mn���K��=�>b~>a���wmA����X>�#H>��C���c=���=9i=�2���'>5�u<��=��$��Y��i>;gѾ�9�=���Z:>\=����s>dӖ=4d>����x�=l�5��q��
U>[�1�7P���M>�3�=B� >vr;���;����>zm�z�	qս`a>Zi� ��J��N4��J	�&��=N�&>媆=MEi�
�>�+e������s�c�>�g��[�="<v=�<G>��~���Q> ξ�E�=c\ ����=Y��=[L����=!]�����=C ?�aBv>�*�-�W�ϳ�G1>�6��7�2>����)��-8�>���>'����`�=p̒>t�n>_{ؾRà��%缏a�=ȗ�>��T�R틾���=��E>Q�/>M�����gc>ӽ&L۽��l�Q>4��G��!��;cm>Y�/� ;���>�C2=gs>��	�'���>�$��命l��;�@>�K#�W'��w ��ۅ�f
2=���͂>~j�$!M�X��=�v8?�p»�
���5>ׅ��a:��e%=�K�="��<���>���^��-��j>k��;�*tX��{>���*U��W���}�>RS\��,�=S��J�>L�%>9/��*K?��<T�s��q>R���Z��=����_ڽ��K�>��>i��F�<lE�=��>��>�5�>���)q9>���=�v����~d�>�!>�����Cr�>D">�NO�K�T�����+�>i�ɽ��@>s��w�x>~\f=�ԇ�}[��>����V��!C��̑>b�4��!�
�)�y��-񆾽�M������s�>��=��c�2M�*n����7>�>��c� ��>�#p>_Q�=�˨�� d����=˰�=��N>������c�,�C>&��>�`�������>�UF:4����lq�q;�=��6>-�?LE��	�N�>~v>�Ԋ�K��6�`�6����s�u�1��!�*<����{*�����O?A�n�J�=i�/?f)L?�X���8?��x?���>��>8!�>3?�U.=�o >��c=��?/*?�?�=�O;��\=N �>��-�zV=\Ď>V,?Y%�>M��2�\c������Z�>mn�>�&�1Cl?�4.>���2->+;�<�ü�t��"h=}4��/�	�%�1<Ro�n]>�־�?z>��=����k=�ʂ=fn�>�W��g@�� ��>�E.?��S�V#9�Y:S�Y��>�E�>���?A������?�d��ʟ�yf_>X�<I��=�����6I�6�s�5A=�i�=�ͪ�WK?FB�> ��=֖?m[ؾ��˾~��>�j�>���=��A���>�]?Q�<89�I4��Q�?�o���Ծ��J�&�k�;6�<�e�?�2���L>^|��A�>�ת��ʾ����>X>:?;����������>��\Qս-��l>���c�g=s�=İ>z��a�޾^p�F��=IП>�0ϻ�$��q���
L����>�����<�r�I>q�U�Ș���4�`�=�b=>i"=p�'�-�`��X��\�3� ?��y���k����=�'N?�3|�7�q�.f ��i)>ڞ߾��Ծ�ⶾ.��>,���鍾X9>��|bǽƲ�>/�n	>��>�Ӿ��Q=��D?nw�>��=3d�>�ξ�T�r�Y�U�&����=�L6��� ���0?<��>	s���ѽ�P�=�E�=�u����㝌��^�r0>!%۾hp?sF�>f�.?��=<.I?o���2��S>&ܾ)*��ik�3�S���#��>�\����0)�>��¾@�!>Moվ�d?�:��
���ŉ<�>)?�q��';�������G>�Nսf_K?Wk>�M?�&���7���Va��Me>`f�>KJl�B����9����1�o���=ob-��v�e��<Q��N-�0:]��34?��f?�5ڽ��9�w?W���LC>�-<m�e>ej�>��>]z��2V���1>�5<��i��d�,?0O��ww��D?~冾�K>Ew�=V��=n�(>6�?��F�[����4�>ע�=; ?TϾ�	?��8�5�Z>'��=.��>�`��s4>Zr?t�\����<��c?ö���L2?���p�C�uϐ>P	��A�?9��<������>�w�>�3���d�� n��n��>^IʾD�>h����/�>�}�>I�ߎ}>iWҽ��z>o�>��?�	����q��>��=�>��Y�?�CF�G�%�3
�3�=	�N3�>3�A��2=�Ã>P*�����?�؂>>��+,>��]�wnپ���=�Y��8 �(���죋��w]>qt=�$��'��%	?*m������9��%B>Z��=B^L?�,�>�d�>��;���m�P�%����?�?���}?�h?�>G>}(����=۱>�^?�����5�9W�?�AP?C7 � ���VG?Lm=
>j<��R���>#Ą>@^2�������={��2���� '�}T�>��ڽs��>'�?nuI�7��>Å[?�W�>�q�>�?�'>��>�?
��=i�.>��O�é4?����+����>4Ɏ�/R�>�b>����q>� �>kv9�7�+�f:>(վ�}Ŝ�Py?Z7?�c��x�d�?��t>�v�=���=T��<�'!>���>C����
?Q09?��a��W��t��4��s?ÛE>@�꾴0־�>�4��ݩ���Ǚ<E�AP>�Q:��1;�}�>#?;Y�=�� ?������>��>�2>��Ǿ��>�Z�>�r?�����¾T�ᾨ�=��7s,�6Nr�
~Y>B�d��S=�d9=B�=�(=]�ͽ�@����>�K�=/X>ٴ�=^=�>>ٓ��B�>��>�B�=?��>>=�:�O>O"h�h�����׍��V1���>��A�ƿ���2�1*>#�<�Rؾ���u;���y�>��r�q��>�s=�i_=�v4>��%>4 U�T��䶡>�)>k*�/���I�	I�>�)����Z���3==�<�l��=TK߽����z�Ƚ� �>�=(�	����>���Aq(>V��>�W޽H���R����?=������>َ�VI'��E���H��}�j\𽰏��C�ڽ�Fd?**��(8��=�F?����$��>��ڽa��=�с�2�`����d�>~Y�>�YܽG{��t#�� �=�ӽf���4T=��_=Y�C� �>���>�['��>ޅ5��]�M��0�G������n�>�ќ>M�>�>�>n���2�v=2�P+&?��G>nRk���0��I�>E�>$3��� >G?�8�>�6�9)��?��>ŬɾsPu��� ���=&����Q�=^����o=�M�������>�M$?��@?4��>��Y>RF� N^>���>�Y�j�J��Z�>�,�>���>��ؾ�쥾�&ɾBB,=oX?�H�>8j?On��Rڽ�?V (>�mI����>��=��?'��<O�
���O����t~�J�����?�8e?*���h9�#�a?��ս��q>�R	���1=} �>��>}�m`>k�=�e>�gE�g�>[6 �D�=4ϥ<٬�=
(�<��=��|�I�Ⱦ���]+���J��n���0ƾvh����Ľ�)�>���M'�>�8�;[0ϼ�i��T?~��>����*����=�P��Q��>��>�>d�^(нP��.BQ>[FL?�~]��r˾����r)?������F,���L�>_F�?Dq�>Q�>���>�|>�?�����;9=	>fj��W���)>����g��gʞ����?��ͻ��-�9��>O��>�%9=� ?DqZ�c�/a
?~��>�mj��1<<vm�>]�>���t�=�'�%���X�q�&������_?���=�=T�>��<����>�&���\����>�?�2��P�����$?>؁?��m?g��>��>���;@o�g�m?E龆�i=>��>F@s?�eм�K��'�=H�����λ����]��?��?i�վ'����?Ad�>��<�'������{>�
�>�aþ�h�>�I:?ݻ�CE>�?��C�8?*0��_l��k#>�(�=����& ���>���=F+���@>����u�i>7/��k?qLN�?�&��>�x�>�ꩿ��潗�;�d���u��Q3��Ƞ	��H�>����z/�A��<���iH��h�>`F���O�e� =�_��֘>�콀��<S�=V�=�������0)?F�����#��G�>A`N�\|~>�O�=��	?e���0\�;�7m>4��=c�-�g� ?�C>�6�>P+-���=�%�f?l">kv�>o0���� ?p۲���<q��\��>���>}��>���8a��2HI<!=�)�>���C>-�°�>�!U>?���y���F����v��8�����������>v+�*�9���=d�3?��0���F�R��>�Z6?���>}��\ֽM�=tR���1��ԛ�[�?����ҿ5�K�=)�|����>������?�ʗ�* ���B>�p7=����쯾h�P9G���+QŽ���>���)7�>er>ݍ�F�n;>y��=^����j05>�7�=�����۾&�a��\�>&�><j4�ck3>jmd?sQ�>�&;>��w?�w�=�U���?P�X>�@���o=�ҍ>�창�+?��нV2 ��s>Ow?���Z��=ޛ�>9�>�.�8�?y�a=�q�>w����> Y���
?DS����`.ž���>��6���l�U�>A�>�UĿ���>i�
���ӽ�����`��nR��7w=�'徛f	��[���$�}���~>�DJ���>ל��������>�$?��=��h�S�>�x�=Ճ�=U�A?2m�8�~�݂c?��PI�>�q��v��:�=��J��'v=���=�bɾ����i�>B��<�O�VY½_Ap=K%@?��=��>��-��?̕ƽ��U�>2����c
�#1���2=E{���ӆ������)>��D>� ?��Z?N�>�2��w@>ǑG?ݰj��C?Fߍ>�c�=��=L�>���>üp��ύ�
Y\>��?�s�>%^���Վ>k��>
����nS?2(a>�U#?L����'�g�%�/th��y��3Y=�j�>��W>�a�?ee1��#�>(� ��ԗ;H�z=�-s>�U�~�V��e4?���>��<%[���9g��}�>�>_�8> f)�C�����~=��8?��^�L�ƽA�h�_!�>��ھ��.>-s�#bm>n?���>VA?[�k?N�־�+?��=;�>Q���?>�4<��B�;G�>�g?ཨ��8�󜜾3i�>�l?��p��%%��z>6��>QM����ѽ�<<>:�?y�;w)�|�p���������N��>�9�Q~��H$=��m��N�v�6�Z���? ?\V2�)�������~ĉ>Q�?x�ؾ��!�T�=䲾g����^>^�T? s�F���4u��6?���>=���4���5
.?�x�=ܠؽU?���'��C^�>
mX�a����?�FӾ�3Z�ң�>J|=
�]>dA�>��m����Q:������>����e��q��*a�=�?_����Q�/I)�0L��K�Ti�� T?�<��S��1�"��>���>�rk?���������E�8:�>�r#�.�	=��B>��?2������nX�J3����s�=�N>�]��T?�t->G}�>��B����=[��=J������5����� ?�s�*s���a�>�@�>�=6}�?�X�?�G�����`Nu>l+���>[��u�W�M���%�>�O�>���@��=�-<�ا��Z�yg�=��Q>";|��'����>�5:>�� �\����>l.?N)�>��I�̕?)Ky�&H���y��ܽa��>`+�=]O:�Q3d?��N>^�ƾ��o���b?�����Ӕ�#�H���K��η>��>-þLѧ�Z����>��Z?��׾��>>�$�>~,?,q�����=��?�\����T����-־�V�UC6�:G-�#"?���	#F���׾/TA?>Bfн�0>z�B=X�ڼ�>v�>C����>�}�<%7^?d��\i�=k!j>�0�=X�`��
��ާ��Y	�D�5�P�`����p�;X?¹��&�H=�c"��^�?�#�u$�<_�>_��>hOt?�Z?�J)?HdZ>��x���K�㽭���D�O�2�>�y?>�J�#��>y�]>2:??'Z+�$h뾬S�>��(����4Z=7�~>>��>hM���G�;OF'�p��>���.�<&,G�=��7�ɽ!bM�P��1����>Ǿ��b�U]�FY4��*�=6q?�M��:�޾	�T?ow�=҃��ľ[�>5�?hi?b3?��>*l׾i6��4���M��k��v��jM
�O��<V���
4?^|o?�ȴ?N�O*�>ez?j	�>��N�?]�?�]ǽ��N��꾍�?~�,?�2�=���4�>�w?(ك�,R�=��?�-,<'`��XN���ݔ�p�?��%�0�Ҿ~"��;>�><J6?q�?)pV�뎟>��R>�������� �=�?{?��0�Uz>������^?4Z?��ݽ��<�Ú�[>�-�>���Si�ʖ�˘a�H����;>�t��a; �$��gar?I�?L-j���}>�	Z>�z�>�TW*?��?�y��>'������1?>�>�%h>O��H �@g>U�&�H,�#Jͽh/?�������v��>Ӕ1>y�>m�b>H�y"?.�>5�Ҿ�)V�Ƣ<?ۻ?���>�락���*���J!o�I�������ڽ�b/�\#�4�>8"��>��B��>�>^�(�?m@?���k����>h<�����Z�> �H�d�>�8*>�& >Rr�e��{)����@�����>��=�0!�=l�?�T�>>����δ��y]��վ ��>�"��Ԥ�]���y�?���>j�&?�.�>#犽0�=yz�>,�2><���D
=+�ھ���F�>�����!�[̳���>0*��h�=-?q�WX�s�=nTj>�=�>zs����#?�<,=�y�^.�:G*?q���Y>���H���9�U�ƽ˾sǂ>�<+��@^>��>�Y���^��
?�h�>ֳ�>^b���w��7�>��[>�+�$R�@��?�pk�q�W�>zS���?r���ﾋ�4<�<��b#;�ӭ�>��?���Bԫ>��ؾN��,ľ��q����Iv@�s�?s��>���ە�>�}b�M����QG>��o��Ȏ<�]۾C�B>$t�=��Ⱦ@�<�ɾ>h�
>

:>=�C=t�}?ƕ�=5�.?���a�>�_p=�����;���c?���<�վ�nx�~�?���v4?zi*?����m�?P�{>ɷ�>��>$�W���>\"���>y�E�)YľP�Ol:��,? a?�W�",?ߞ$?�ҥ>�6���<�`+?����魾=�=P��.����̾Т�s>8��>+���d�侩����>"�Z?���Z3��y�>��,?���V�+>	P?1	)�/Hk<K>���~���gs��>��?�Tb?o�)��������5	�d��>�٣>K�55��(�>lL�=/pw��g�>���m���Ӥk>*��IڽI�A��x1��}�>>9,����=A��>}�6?t$.�����^>$'��QA>���>E='=6A�����̬��r^����'?��b?;�w>~k�>�\?�"�= ��?F�?��k>����>�p��P¶>�0T��������������5>��>U�$>�h<>�U�>���> �s��&�<���>:8>Hۺ�1~>:�>@f˾���gt�<��<���	��HA���c��[?��*?	9>�������%>=[�?�ʴ������Y�=����ܺ2�5��>|��>�	S�۟>�����IH>�>�� �4�?bRR=�'?8�??��b��)R?Ȭ����R��:=�_��Dǽf.�������ki>r�徃��o���-��?���>�x��L��=ދ>}q\?b���.?yÀ?'k�����4�r8�>���9m��8n���7?cQY���=@�>�>g>��d>�Ԛ�y0S=��w>�Ǿ�Ľ
L�>�z��*E?+�!>���>8H9�-����!>�L��^�����D��)?_�־�u���1<��xվɝA��'����=�E���,���>�U	�Q>ف
>��?�����e-��>�>�׽G u���ݾla������8�>5/5�CL�?�@=R#>���>n��>r|]>7o>71�>��>N~O�-9��uc��i��?��B>T���ū�����>OFU?��,�䰈=�d/?�f>�n����T�3�99S���$=��g>3����>%��=�q�><le���� >Yci�0u{�:�A��`�>�,�/F��04$>�^�=jo�>��>�f�>�oڽ9_-?M/V�Z
���C���j��ɯ�7k\�:33?'n꾝ֿ-�5��ص�Ѧ�<� ���?��k��>J�?�.*��+�� ?���>/NB?g�E?~�?��S>'��=]K�\����X�=�?3�<,ޏ�r����>26{�H���Z�轥�_?B����Ͼ�?�X�>�-�=��s?��?���=#h�>�Z��!��*Y?���\��<$zm��<�
K>L�J������G�֖V?��T?`�>#x> �?�9��v���?���>�R:�Շ�����>6&�5�[��<�>#f�|�/=q��j>��ֽy��>��x_�Wm>�a���	�!!9����?v쀾זi��>ڽw9� �8��p���=ɫ�>�	8�sžrCy���?�CK?��<�z(?����oV�=VsM�8G�l�ᾄ.?_�?�%��9�
��h�	N	?'���������y��6i>g@��b�&�"�)Iľ���l>N�>�>��H?�+>�K�<����=���f�����iJe�ݚ.��Dս�K���⾩1�=[>1u�>�i�?[K?6�<t�>ʆ�=R��?��=�>`��>��<?�f?9�>��>_�(?'>L�=�a1?���>��չ4>yJ>��X�?w	?���>%ى>3܀��sN��Rn�_
��&Ƚ��?-��=�%�?�-�>���>�b=� ؽ�(>Q��=ݞ�=	�)��RI�@J޾�H����"?��5H/?��������G�w3>��>?�>a���
������=�b����P?��N?f�D���=�W�>�[n>���?||�>��?4-K>���>#>�f����>�U7��6��*R>U������>�]�� m���hj?��$<���>�>�>G��> ���e��>*�_?�Q�>7\(����>�R�ξ<]"��1���>��A�l�_��Y�$�5�	��>�l�>7�F>ۛ��C��㾠%	?|��?-��=ڦ/?FV��ȩѾ_����� =+
?r�U<:�>=�T���?����(��=r!��U�>���<-���E� ��>�O��c,	?�Rڿpo<��z�&t���a�3Ͼ#o��I��G�-�Dl���
��>���t���Tf�� �K��x/�:S&�'����=a��c�=s.���ؾU�;��*w?�"�<��R)�>�l>U
|= b?L�辕�/>����zW?��/?$�v>Y��>���<����)���D�>^��+����b�>6#�d��?����K�=���z�<Zw��C���/{о���w>u�>
+>w	�>���>~'�>f,�>P�?\ӻ> �N=�����(�[��>�f=�}�=��/�����H�o������=�={>����*�t>�Z�>6=�ᬽ�6�>����)	�"֩��g>l$�>.�c? ��>z�>�s���>�
����>R ��ڴ=˞?$9�G���&=�ja��o����>A ��z��I��>�����
>i�g?(q���h��W<;>~��;_9>�ƪ����>���>�"�>��,�V�оrD�>/����>���=���R��n��,�<�ƾ ���iv�UE"���o�^'�=锼��>3�?��G�	�>�� >�.�?�Md���>�AO�ҽ>.X�6}����?ê���g�ܴ�����E><ؾ�j5���=91w��^�?\~�<�8�<���=o�>q�����޾ P���
�>k٦>�(�?�C�>���>�5����X=1��?F�X��L��Z�V�t�?�F&�Ke?�4?�%d?㸵��i���n��k�v/����=+�4�:LP?�a��X!U;j��Ի�KT���"�>��3�YfR��0��{,�f۾�ë>΄�5�>��&>É�;�����	�����4$?�k��/,���%�X�?	�>�2$?��@?g_?��)��8���Ш�2�
���վf��=�������?�G�>5z=��=�a?��*?DO�>�Z.?�އ�!��>���>��?t��ĵ_���>4r���<�>�I�=��$?<n�>�`?K��e#?3+?\�b���u��&�=d�>f&�_z���:��D9�>��>#>o��>o��>$&?�t >'���H�?1��>v��>í->_�>�ą��^�>gW?�Ҩ>��=yAy����>�T6����D)Y>����� 1?OW����=�JR����>C�Žr !>#�>-�$>��>�\>�+?�ޮ>���>B��r�?�}Y?T�=�j_=���>}����>��𽂌�=z�u�=Ju�d��������<(@�>�Y��Ԏ�~l�>$��=Yu��ƝK?\F]��p>�L�>�b��&�����	>o� ?u0?>z;5��x<�P�!������1%��B�'��p���L��0������<����YbE=��e<��>D��>�|	?�2�>'��>��,�!�>";� ?-Z;��������薾�Ͼ�J��(1P��#>_���=�`*��ꍐ>|�쾴�"�E�D�
@�R�/=Z��='5�>���< N8�(q�>y#>�Jؼs(>���>5`;� ����	=���x���v�ￋ�վ��#���������g�kU�����>q�>���^�$?R���>���J=�K�<'��;�K�>-A����>��>�j=�ra�N�=K������M�ۆH��V>�>+�Z��?gW�>q��=9r>d����F?���x�O���B�\"�>���:��$����&��TO�qc�����瀉����=b:���d�>��Y�����=ľ騖����=�9��q�Iv¾hG��O�>�9B=�B)?Ͳo>�Z�����?������5z��?��
��7��M�>���>�.=%�?�!̽��?���;��1>�ڹ��!��2��������}fI���>�5ʾ�S'��W?أ�>~J?5j˽�a�>�-�>��?�`�=6�$>�Ӿ(a;�\N�r��ء��{�q�鷈���l����˧�>Ic�?tK?��:?�?��.��#�B�<�Q�>cv�<'�)���Z�F�,�ze��6��
;����{>C�^>
�=I�f߮>�o%����>&ڃ���>>��>�Z�>��<�hJ?y��>l�/=�����>�4M�(��>����vj>m8?|P?�����'�08��1���w9>�,�>�n�>TK>��>�h4����C�r?�z�=�a��/�ϭ+?J_{���a�@��F��>�Ի>M��>ϯ~>���>G�>�m>h���e[�>�}�=̌;���9=�WI>q��=��cAJ��t�<�?� A?�0>�6�>��?]jt����?rj�>>s㣽&h�~Q_<1c(?�n{>͑���>g������;�>�~>��>==��>U����8?� ?�X��E|)��Y?>�ʸ�V)��?̾@��|q�@�8���侦)<��?'P>�>}���y%>��7�gݧ>ߐ�))"��#���^(>2c�n�J?�yU?��<��>)#?i���̿&?L��>O��>;�5?��>�?�L#>�C�>R]��>�0>�����(	�=l+;���=έ)�σt>cT&=�r�>��>���=��>²�>M�>�Ī>+�|?cN?^D����1�H�~��?'�����=g�@��y?���O��<뺒>d>y(&������p����7�Q�cF�=G�?�Ծ�s�>��<a�C����,�����<�����o�C'�<�>};}�C�+�k��<b_�:�I�2Eɾv(¿㾴ʾ.	���~�>J
$����'�6�M*�>�[�=nw&��>�6��֔==�>��M�>�����s>[-�<0�>?O��5`�>ē�>F�$?�����+?>S���U�h��(׾�"�=�r9<O9y?!��>S���=,���L�=B�8_�>�i�>
��=�龺T���M�>���=��.��_�>�<�B��=�瞾������&Wؾ�0Խ|q��Іݾ!���ĉ��-v� �����<�P���d�=b�����>�ǳ=ӽ�"�>Su�L����<�/?�&wC��ZV>�N���Le���Ľ��پ��'=��0��x�?F�ǽ ���Ҵ�>�1%�\j,�L�ܾ8.
=�;���=��>U����?���GǾ�M�ׅ����>m���W���x�<��о&��Qf%���=W}�>f1�=3䜾��=>�F�>��`>��4?�.�?�Z�?��(>0g�>�����?�]�=pP�>'�����$�i��վ�eB>��e>�E9>�*?��>�a�>�?�<kn�&�Y.?ѭ��$��yq���V��e��)޾���=Y�F�g�>i؎���T>���=U<_�cXF>�4���}��D�=գ��"^����>���J�3��y6>WA�(��c�>&[ ��$��G��]M;��׽�;�=�&�>��?�@?���t	��%?�Oڼu@`>p>g-?�3;�"Ć>�ؾs{>�{v��>>'�ɾ؟��>��`/��(<�Ȗ��S>��[?���>@|{>]"����s?U�Ѿ�|8>7�ÿ�̽�8��Ā�2R0>�\>�&����GSv��q>�T?�A=��T>&���:?��>1��=��^�\��h`?�	�?��h<_��$i��r?}W�T	q��<�J>��	?��=̡�>tZ�KG	��L��S�>��~>��A�%G8���S�g����&ܽM�7�WT�>G�9?Г�>����I}���(�J]�R�ӽ]��.�?��]�/�
�y �_0�>EF$�i�>?��>�Z�?v$Ͼ�<�tی�S�n?~-?'�?�~>��G�hk�Ņ�<�?/�>kЋ��n$?���>f,?ȴ羴��Bľ�ϩ>7G2�����א1�)��?d��d�B;04�<o�>H���Vd�q?��1>�T�.��=��O���G�ep#�-!�>��>?1�=�A���\ۼ����,XX�R�,>���0z��Q�b���"?%�2�x	�=I�ʼ-Q(?���?����e�� +�I;�>�4l>�ݛ?��?������M=<���F7?�I���<Ta�=tH�H��z%x�І�ѫX?��;��=��x�>>QѾ,���H�;�a��]<Ӝ�=p��>T�.��H�>�j�?^=>���<�L��H�G�l�?*j\>�@������;?8)�/ٽ������>Ģ`�PT^�Gm�bU=?�A��3�6W>{۾��?������&�9�Ǿo)�>�����^�;�?�<�B.?a6�?�Ŏ=�оU�Y�������9} ����ÕD��n?�\>��O`�=���>��ѽt+Ծ��˾�D?�O	�L����>�� �>���>�?�A ?2��>�>�*��?��>�K:�AT�vh��^��9�0>
�q�_^�56$=o��V;?F �)Y�AV5?hq�>>�e��=�&�P?v��>>������nD�k�>&?/ �>��G?�n:�|��K1?HU>׳�>�R�>g�>�F׾� _�[8�=�?)�}�Ln�Jd��n��~�=M�<C�?ޢ{>�?�$�O7?�K=飞�pQ����-�^A�?hm�=�{��S�>:�3�so�=`�x������������g�����������?aB?3��P�?�F@��t��=?$@g��?&��>:@? ii�~g���Ϯ��;?���>�/H��0�~�=��?������7��Tѽ:|��/iL�#�P�˓�=���?!H>��{
��=.��>�����q>贝��QC?7=�W?�\�?��?D5>��=҅M?Z���W�=5�+?��0?�����P��Q�=�
.?�v>n ����g��M�zp��?�u�2��X�˼�<��f7�g��>�J�>u�M?�x'�pk=��V��LG>��s���2?p(3��K�����>��7=�J�������>;��>�������C5�3�	?�W8?6B�>�e�>�@3�i��q��� x��t
O��J8=��5����>6���3�k�=K��=N*?���>X'���u?}�D�ti�<z�+?�?�b@��O>��4�k�?�s��?��A? �U=��Z����=��;���=+?��� )���	2�.��>��?�	*?ˆ��KZl=��>??�>��C?���=M]
?*��~OB?Қ�˷>�@�%h?�,�K	4>{�s�%;?�	I?��˽�>6>�KR�Dב> �B��z�>.�о�ͧ�t+�iS�>��^-���[�>��ľ��>��"�Ң&?��>���oo=���#=?���\66?���*3��Ss>Pb-?�LS���><����\+>�VU�Q���C�d?�>�֩���=���>:�>�V�?\�o�z�6����>巧���c?E�n�� ���J�=9�E?�f>,|e>R���O`���
F�TD>ZȒ�� � ����=�A
?��>�پn��;�?��>Q�b�!o(>N�L>�c>7���v�#j���ҥ>�Wb=��E�ك�>(��:(}?��h�ǎo��A�>:���X�>����r�>|ў=����,�><nS��t�>����A&?�Aʽ�J�:���S�?�nZ��/=�j2H��I��e]�ލ�>���J�!�ij%���T>�"�>�
�>�;9�A}	>~��>���>�O���=�s0=v,T�����^���՝>8bP>s?��?gh�����]?�����| ����M��1N��?*I�ek�>�(��u�<���y�=m�I���?���7�0?*N��\>9����a'���4>��B?EA-��]8�\`	�fl��%�;�d�����ަ�3v>���>�~�>�@���P?!�]?=*���<N�ξug�tk>˂�>�>��F;�[�>�l��A���q��W?��}��RB�3��\�>tl�����>���"��>\��=f)�;�*�=R�A>ήļ�1��p>jz�9M>-��g�Ra�>퓧���i�w���?lk����a?�>Z?�b?����G��>�9Ծ��5?��=�,��[߉> ���M@����2�����%��=}g?�!�?D��}�t�����v�B���[�Ps=с���>�-?��>��n��h�
���ݦ����,?��>��>�链��0?~��Y��>Y[���6g?�T$?��֐�?�#?$�?J�(?2�n����7�?T1"?������$���V_�?���;�?%/�",�����Ǿݻ�>M��>Qv�P���:�Y�Q>b���	ݾn��/u?o?B��o��;��/�O��>���iw�?�8$�i�b=�'���W!�=��������>��> O!�Ԉl�*�׾���>�O���b? �o?� ?!=�?��=��=�K�P1�>�K�zV���P�>R{��=wL�߬>��?�o�dS�>&C����>��ѽ� \?�����_=��0;����(>��=���x�=
 �^���{C��T>Uz��k{���#?gN>���?��:=Nt
>9�6�drg� ��=��m?f�>(��>VJ�U�޽Վ>�R?����s#�>�>#C'?�H/���=�
��>�| =X���A�{?6�>�׾m�7��4�k��g�������.��!2@>��;*ӕ��	{>���a���Y��]?S�	�+?�ްO�/Ƹ>9�z?�> ]�<�D?��.?Ն�����n.?��K�7 ˾�����>��?�m�U}�=�ʴ=���>>���n�b?%V�>�p潨^�>��?K�Z�r��>�+�Vڵ>1$-�[/���N?�?T�!��j��r�n��=*p�$8Ǿ�¾����v�>C�2?j�$>qr�=y�>��?��D��_��jn>n�ݾxQ�>�>��>��>���th߾m$7?b��>x�2��0���=�l�>�>}��> 42?�D������ړM?�4����C�^%�]Ǟ>�~(>t�6�pj���e?�e:?�P?VH0�a���gl>w�3>��?m >�s��?M�R��?<�ؾ��>������>Я����;Ў<?��>'>ͼ�O/�a���=0?�L?��L>"��=isq?4�-��>��}9[??�(��Uþ�=�>�)`?T���%̾ 3Q�Ġ-���v����<��?�&�=k]m��^�>S�S>0U��t>
�&��-��#���o�<񯀽��B?wu?�3�1*����'�>k��=v�>U��>%a�>�(��Vk�W�>��?qJ�=&�>����UV?e\�>w�˻�~=?z�?Q���!�>Y�k=+jμZ�7�����	�>�I?�~��a>�4�
��?}�4?27���UZ�4�?�� �x�9?>��Z�>�s�;�?j8J?^�a?�����+����@��>)�����о>�,?&*����>�O�t��>�Vھ���ܟ�\�>*���Q<��z3��?f[��h+п��J���?ƅ	=���<�B����D=�J>��?��>{e�?����.��B�?�ؒ�%��?��i>o�>c��=꼵>�P��*����g>�	:?�.�8Ï�����^=��W?O�S��:p=+����[=�}���]e�M��h�v�fD����<==y�����>�J
��\ҽ����N����h+��=�̠<߫3=H�k<�Ȟ<G�<��Q=X]��O�J<Dq=��l=NX�<���=�*�=�,�=l�$��z�/l=�П<���� ��=�Y<�Ɓ<��4:��;��<�"=��m��9��h/&��k��U=߃�=��u=U��=Z)=���c<�U�<p��<�̄<;´;9u�<`ȑ=��'<�ͮ<�=:�=��K=��g��:=�,��7�4)�;�==g��>��<����X�<4B=T/Ks��=b9^=�|�=㵈=	Me=4��<�AW���=A0�<r�;�}:�����=�u
=�ϼ��=�Y�=~�,��~<$��;�3o�;�$�fEg�d��vK��cĘ��3�<�Q=���<s3���K��6����T��m��=�=&<����R���0=��)�d�K���Z�E�=��?=��:7����k3<O�2=���<�HG<Y\�<N���돽A��t+M=(S�����rٵ�&��<Y}�{&��'7Q�2wh��)��4�<W~��P���3�C�߳��7>K�F�S��I!�ȡ�;	jԼ>��"�̼�CP��"��X��+����M�uWJ�T=�a�	�Y��hc�ꂽm�B���ҽ�߇���?<�I���m��kㆽ�Q���Q����Dݿ��0����<��2�~�"�?�բ'= V�<ex)<�P	��|���	λB�<�u�𶞼H(��'����<!=�j�
=�'k=3=o�3<�;������o=-ڢ���5�s�c�^��=#D�;'�;W�k=��=�Ğ=~ʻ=*�S=��;�����==y�=�w= �]<k!����<�~�<�b���ɼ��:.�=۩��")b;�{=��<.�<e���<9�u=z��џ�,(=��=�3=�ݗ=�@�=H,=�W*<-=S=+"<�GY=��C�i�1<ɵ��'r=����󏼊xl�4�]cu�%��BX}�3L��t<Z��=Kf�=yb��;�=n��;�A�=ND�U07=��=���=�V�<�_>=8ţ=���<��Ǽ�3�1B������˼����r
��7�'���x���3�P�C��<E8��.J=����KT�<�m.<p��;�!��dz�c�<��C=�|<�-��\=�U<�:������#w���Ň�
0�<VԾ���:��=G<��g=E_�Io;�[��+=X�,=����:�;=
R=$q=5[�=V�=��ͼ錠��L�<����%�=�E�=K{�<��Żm˧<��;��_=}�X<�f<�3_=��<A�;��C��@$��FD<{~���#�_)N=>b#=� Q���:��I�<�T<t�b����^:<6���f����6=�:���
�<�L;DӺ�&��
T��E=��|<�,�;~�2<���<�
�=��O<��d=A}�=3^g�;@=���������<̝=���43�=ܬ��F#o=���<y��<C�=���=�O�=��<��<��R=��c=`\�=��z�)�5=�-=��U=|�����<'#&=r�=�*�5=�^=�x=˼_�uNA���e=�lS=.v�<V�9=��@<]�=��$���3=_	Q��P=�m�=�*�=�:J:�;�eD<�/�=�N�=꧄=�|X=��:=��<���=e��<H(�<�>l=��<=Z�_=l�e�}oܼ��9�d�<5rC=p��=;ي=��H<MT�=*��=e�h=��&��o=��=8<��&=�Fa=���=�9.=7�<0�<͠=��<,��=���=��-�<ɵ=�;ɼ֪K�� �<�';=A¯;��N�B�Ȼ��*��xC�h^��*��Z\�<�߼6���N�[����	g�_�;��#����	-4����]�Uw�ĉ��f��K���
�a+M=��+��l��x���<F�<������7[�<�I �%�}<1�j�S�%�l��1!S�ᘽ)���C�;W3��ռ�l��X*	�!���J�=�}=��oj�<i�=C=?���P=M˼�V�<B����=B�<�sh=Ùd<d\�<I=$L�<�|=��?�	_d�}">�"�?�� ���(=l5�<	��b�;;���<X��<uBn���I��\K<y��<1r���������qܻz�hE�<��o<УL�JAػ�,w�l9 �G���i����/��č�ed����=1�+:;e=�Z}�} �=G�B=E�K<����*g�=�ǡ�!���i�4�=�QU<Y���⳼4C���rʻ|
	�YQ.<�����𞼳�����R��hu��� :߃����?�ď������d�;�7���7<H(�< ��<	3�=[�~=�;�C9ȼf�=��F<���:�ۼ#� =q�"=�P< d��w��<��=B����W�4�=�u��P���$�9�́= U=}���U�����<�L=���<�E�;iN=�<$=v�\=Y�=���=��h��NI=�S=�*~=���'������<�]�;Г&��K<��Z�
۱�O����ù��#;;{q����>=�m���S(�����ĿǼV1�;�,=�^���O���s�`:�����<�ip=OF�=8��=Ϯ�z7^=)��=Ξ�=)��<���=�q=�R�==Ǎ<�j=,P8=�ت=�=�T;=��%=٪;u@�<���ux�<oԬ=2@7;� �<�����&��+d�<J�����<׆9=�z�<X�Z;_� =�a����h;��,� =�2;=.F伄ȯ���<�\�=>��<����Lu�=�W<0�L�JV��ʉ���z�.����0v<W{��dY�kBS��h�����=��5�n��<L�=Z���=5B�<Vk�< �	=���;x��=b��;��2=#^=GK=J�*����< q0<�<ڀ�;a�];�伄��;������z�<h�l���-���[�;���;�t������4�4Ͻ#	���f�=�D&=��<�����$��0	���=�?ƽ��ʼ��i=��r�_���vG��6��K&�={)#�w�m=]�=s|=��2;V�=
F�<��==+�Q��=��<�֋=u�j�ݦ�<��;�2�9v�'=�=�=��=5��-��=U�s=�@�=V�<䢶=y��=nQ�<6�<";�=/A=�=������s<I޼�׼�㿽�<�8=3l���F����;Yc<;B��H\��)��<�Q<Ϛ�?�$=+΃�<�0<~���B;��G��	�L<�`��n�;��м*��+� `̻вO<�AD�^6d�f���:���͉��/��Sd1��U<Y�1�3���CN#������;�8��f�J�x�<݉\����H�ȼ+v�����j���C1���=�,=x�.��bչ�f!;��/�E�w0�O��<��#=����R���G��=��=A2Y=�X+=s�C=	y�=6%�=�F�;���<�ݭ=��A=��:W�<�Ȩ=���=�҄a��^���������(�L#W��_k�G2��â�}㭽�j��%C��L����v��gvT��(�˛\��`��ꝁ��N�<��Ž�R���R�E�<t��~���_���a伔������CbS��x;��&<�@
=�k�=m��;�����t�8�=Tn8����<>��x�F=�F��6���@��u�=���<zw�;�T�<ȁ_�[Th=T��L�;��N�P;�2>�	;��V;�xy=���+��<��=���<"@J�
��<��k=�l4=^8�<��O=ҷ�<o*�<ؒ�<��<��g=Q�7=)�u<�h�<&�<f`�;_.�<j�=�q�<N��=�A<Qf�;R�����=/9;J2<�e� V=H����C��ݽp=%�ۼc��VN��0/�HW�p��񭽱<\<I(��ߏ��b���V닽m���&�T�3����<�_Ƽ�;=:�6U=���]�=݈�<�$=��<��<=Q<$j=Lm/=��w;U=&=h���t.;��3�;�i�8�<{�ܼ����@���I<�h��j��<Ù�/���0Y���<�>�n�=��A��;(>��>��
�h��=�Ҿ=�"?���%�'�"�)�aX�>d�4�v�߽)r�*�G�]���J�>˅D?*���͂R?>�Y���(�>0��|V?��?���?�W>��9=���?홱�%y4?��=f"%?��?���>G�F<�N5>�Y��|;%?9�>��>��Ҿ\�[��7#�=ր���S>��
>q�>�/%?�g�>�W���>q>������?]S��L�59�=u&?1��=��=�d�� ?���>1|B?�QJ?��l�������~?�Gi��Lw>lG���<=i�����{ջǭ���i�>.��>�:�>�|*?���>�
���m?�IC�*�?���aS��G]> �1>W		>����?��w��ߜ>3ڼ�>��J>���>_�����r>��,3?���>����ؾ�x*���<���t��<��н\��N7�D�@=��B�UQ����"F�>��=ͽ��z�׾i�?��^��['?���>�4;?e�?V��<��B�re>>��k��9��ڭ=��>S���۲N��þ�\>��b=��>|�=Ɠܻ�ýN�Ծ>�%�,�?�L�w��0��=�Uw��59?��콗�ھ��7���۾�n�=�[ܾ e?�%�(s��}8���<��=��Xļ�w�-?Ct@�
B���E�?ϝѾ̪^>��s��h�=[��B�>N�K>��>?m��>�a#���
����>C�>�?vC۾Ͼ��Q�1��+-��u�;� �>��:�>[j�=�5���=߽z�T�0��>��Ⱦ����K�>"��>�=(�XȰ��0>Ο>��>���>�3?{� ?����lW�<_�o�� �>_�,>9�������:�r���f��<�i$�]_��Kg>fT�K����rY��lN�=�>�?h�����2���?=[Di>v��<��>=�>8}S>�Ϲ�H>�_?1Ǵ��Uy=���=
������>,v>�>�E�>LM���j�>޶�� r��H$N�0�B���?���>������>�Qڼ�;�<�ۨ�<ё?�!�=V/��Y�=+Q���+4>�B�N���C�=�M>�&���9>��az�>:��ߊ�3��>���ቿW	ؽC�>��e>��>b�<ք����Ⱦ_Sļ-�r?�e3>��,���J���><[ ? ���W>����l7e>�r�����SH4>'RF���?0P�=8�����>�L5?�xI>�ET��0�J?^|�=^�>��lF.>4���6l2�3���C���s�(>
��>@??��������9�>+v>M}j>67>�d}>yT�=Ⱦ�ԛ<�Â�W�>  �}��>���=1D��o����U=��>Rx�>эV�y�l��L�'ݣ��W�~X�t�~=���=����<½��K��=`��>�̆����6L����=��>u*q>��?fS?D{<T����Ծ4�2�j7���خ<��">a� >#`N�ŕT?��>?�e�=>� ���?N�	�?y�>�2?/u>ǉ�)ձ>DG�<n.�?����m�>h��>�T��7ܾ�>j�;թ?g�����R�w����J�6�]<C?C��	Z��A���w����?S_+?A?�C�><tZ>�fE?;p$?�g�=��?�?�]�=��)?�fH�'U(?@�>����?q�"�W�Y����z�Ӿ�A�W��>�g�>@�U={���@A�>8�<�(�?�)־x�?�M�>`�>����:=?}A�>���>���j��k��Lk>�Hy�����L�������>J�q�I+��kq>���>7�9����X>4�=�!? �>c���>�V�=D>�����ؼ�^?v��?~5�,�Ͻ�����j���#� ����o�p��WT��վ禕>�D���*��:�\fJ>��:?~�=j��=z >��>��=�R>V�#��;�IL>�AB��X&��5Z�9)�>SG=c#���t��q�?�� o�>?j���H>XȾ��[�微C�[���*)��t.��h��о'�"?'XA?�p��$2���m3?�>[>p8ξم����ᾓ�G������/>p徧�>�c�O$�=�#Z?�ӽX�w��v��C�=A~�>r�x>��]?�s���̾��?~L����t21?���=L�? ���'V��Ͼ����Wt=�ڽT�7?��Y>�f�#+��h,?��A��^�=��=�è>e�>ʹ�2z�<��>��`�>�S�d�%>o2��e���%>�`e�鷌<Z�U���>�&��Y�e>�q��r�#p����j<C��F�=�u=��>|HP>�|�>��0�¶־Ug�>�.{>2a��z�侖x���>f�Y�U�ľI'�>��>*գ=>s�=��?��=�Ⱦ��=ʥ���&9?[�*�
��۪>��>B��=��Z��P�=s��>�?>��>��Z?��\>�%�>�q�b�t?�Բ��@>{=���P>C\��#�����m8���=�D?�>�>c�)>��J��?�Ы=X�Ԡ����'=;`?#�	��\۾'�J�0�,�O���\�����>b��>|�=윾��>T��<��>E����;<�>TC��0v�2?�4�<8��>«�=��>�Ob>�,?�^��C,��"=(�>��>��J��y��Ў>�����>�o��Dv��$�=ɝ<@>򰠽}�=�(�O�E���?��+?��B���	�2�m=��c>�'<����>�:�>s����B>@�����>�� ��q(>���S�X?׾���$�����>��=[��>wm�>0H��v|B?2l�>gk���\�?�ɾ�+���v>���>��O?'�5�J=߾��?�!��C��H(>(�;=d?�Z�>'�&�D�?���;ȯi���2>��.�!?M!=p��.EM�[}��_L�<��A��%�ޜ�>��-?�b?1�K�{#�U,�=GXF?���y��>�亽�ް=ԭ��˾�%I����=y� ���?.��;ѯ'?���>8B>s�>,�=��/>�K�?��M�A���3��9mK<�)�>Fx5��B����}>Ѫ�>mC��	����<w=�=8~?-��'?
^j>��<�Ǿ��=?��?��>��>���(:�;ޖ�=ż6����?j�+��u[�=8���L>d[?������*U>Kn>?�X��=�0Ⱦ�^�����=��b>_�	�d�*�v[G��t?�6�(����ry>��T�w���K�վFc"��42��`������͠���#?^��sl<=����%3�=�}�?�$�=�����)>��v>�_�>�1 >�^��Ž�t��^9׾��;?S�?�>	��߬�$?�>*�c?h]={�Z;�?� �>.�~�����I˾e|�>þ?H�>��E?4�==�}����A�>ʉ�=2Qq>ڽb�=g%�Y{�����+�� �̾�?�<��>'���C��a"����>���a���B�ļ9'�>5�N����fР�gx�=. ��>W����P>ܯ�>����TW�=��N�@O?�$���88��q�>TJ�A#��<W������׽��>Ur?��w��*ɾֵ=�?��B�?��N����?CLo>BL�>�f�<� <�
d>���=g�¾�[?����<���T�`=q��aB>z��KH4�&����\�>���� �=~X�>�cm;?���>,1>;(7?�2=�#�>�R�>�/�>5��>.�
�5D�^�,>����0�i=�is��i'>MĖ��ư��>!=?|y!=BZ>8�0���R>���>�$�=�����?
�~�e���~�לq>�ľ�F�Չ�=���L�
���=E�;Я'?����s���=��=��G�3�M;����^V��~�+��S����ʾ2Cy=`�Լ����s��z�<���>CSx?���?o�VaF>�f	?��Ⱦ���>��?o�@=Q���v��?�w+�MV?~%)>X���ny�,4½\㋾d��\$����?�׾Rk��:>@��=�ې��Ō�i�N>�>�>�c��\N�A+Ӿ��(?����� �����I?� ¾%�����>U��?t��>)�<��=��(?��->�}h>h�=ּ*?�(?i�b�F2k��6����=�de>TԠ���>��\?4�?��~�Ĉ�>��u?���=��.���Ⱦ���e��l	��r��?���9�_3�F�>����s�g��D���B�>0 ��������������h?����{"�<?�]�z]X>ʸ�=X�i=�o����>��>�@>~J�����U�>��1?H��ٯ����>���>���?TJ_?(�=�@>��>��̽�j]=���>����/�=���>\���\�>2Nľ�خ�$��=�`	��2�=1m�>,H���� �P�"?l�?r+�� E�>p�>B2���"��i޾N�<A>�	��Y�t9��2�	��9>p�\?�[ѾNgF�z�-=�L�䩾c��%�u���s?��V>�
���v��t?�S�=k:>;Ev>�8>>�U��xO��ڹ�W�>��a���6�	���v?Kr�aH˼F������&��
ْ>p���<��-�>�P�>�*��6�>归���̾�䀽3)"�E��h��;�)��2?����B־�w�=�.?P)��bC���=����V�W����d�b�??�tZ��w��I{�v�`���߽T�>���j�P>��?3��>�ד�d?<�VH=�W��17��Pr
���N��%ڽ�u�r
?D�������>�S�>0���0�>k�Y<
!�>x��zv�����Y�>(3����>��C>��T?L;�>�X5>�[�>¼A����n�>߿�>="%�+�1=M��>k|n��vT>�=@�
�Ҿ�DS>���>L�� (����>��̽�vH�[�ӊ�>���Pܾ]�R>�q�>	7�>��1=�d>�c�>O=���~��.�'>�B�>�/S�IS6���=�>;���o��(ľY��]8�<��A����=ޙ����>H�=�]E,�$�,�y;?�K�>�м����8�>v�!?m��>��D��R�>P�>/�>�� i�����&��&���݊�>< u=���>�e���D��>�豈?�O��8�>j+R>^?8»>��$�b	>;i޾�M.>�J&>I��������>���>2�����<�#DS�<��-�!��;Ͼ�l=ἅ>q���j��>���?�m�ZHx>6j?��@���A>8��>��>X���N<?�?"j�g��>��¢���~���Is�i]>K�����n��=��?�P�L����_��; �=ٛ�:�����m���<��\>z���/>BG?�w?�%4��eV�������lP>\2ս�H�l�=,dc>���ϳ>������=Z�>@f�= �?�k���C>C5���ľTq;�A�>��>��w>���>z�>NӾ�.>�䔽�c��#i?���>M*[��e����>��<����+q^��\'>+tN?�g�>.���r�n)�?���>>Ž��<o?�s>0cýF}¾��<a��>ʽ�>��Y�8ǐ?�(!?���>'�r���y���Ǿ�8>i�<S��>"�*kҽ<i>�ϛ=e�=�Kr>&��>p��?]&v=��?��E3�T�/>�"�>�e�=:l��-d�>6�>��x�V��>�/C����>��=�8:��� ��}=���>4���U��?5�?�LN���$��!�?`׊����Nu>��D?t�4>M����L?] C>�e��[?�JD���]�>�1�>�65��蚽���=D,�>����@ �:!�o�>0 �2N�K��=TB���z���(a��8��ι>��>���>������2?ٳ�=:˾E=��k&R�!���A�������^Or������I�ݾ���]>��o��k����=���=jq�� &�>9���b��>s>�^���?�k<!@>�ʛ>�\��`�Ӿ��1�J��>}���Ezx<��'>x��>.���$+C>@�J=;��>`%Q�����b��ć�t�>��\��`��jƭ�X�ѽO�b�Yޤ�{�>��V>K�!?{Z����Ͼ�w��<�+��Ԛ<\�,���l>�l�>.�;�:K���v�=����jǾ���>��7���>M��>��Ὡ@>?���?D!�>u�=M-�=@ei���"�|�v��μ��𾧃3��U�����1��Ԇw��H�j��?�P-�2<-=��#>�F`?�����}���<�^�>�۽�E��q�����(?a��N�~�Y�������q	���L���#��M>1v�.J��k.���7�ڛ���*>"�����0�@��+g��U?X�<�ar=�;+?�1ľ-P���(�<W�~>��>��b��qY>��1>�e�=����w}>!�>sxY?ں>��O�����>���](�"�:�49>�s�>AOT�gX���qB�5�>�x���ώ������+�B>b��1<W�D���*�1?W�i>Q5P�K�v>Z�Ƚ/y>�R ���m��L??��I�U�4��<���>�7/?O��>=�>�y���y?Wd>M��������o�Q��gk���.�����?OC?�W�U��m�?�	�=�ˢ�ef���<Q5q?�@�>�s��M�L?�wM?E�S=m�v�D���@^ <�%�V��=����`P�9�4j�O��=������i�U�D>|۾Y>�S��id�-#D>�Bx>qy��?�>�1�_����u>_{�f%	�@"0;a�u>:��=��o�^s>`oQ>�5�>l�>g\p��D3>���>����s�U�>�A���$Y� �>8��>-�
?��">��r>|�?=�w?���>u�>��>4��(�3?)>?
0=?�v>�>�͐��Ry��m?ejU�Do�=��+��P��p��ϩ>��I�$C��5��>\�>�v����>@|�qR�=#:��5�����3���'�<R"�96?�3>��>�D��\�>��e>�=:jv�9U���?��?��I�J�e> q?��>xd,���0>��=g�	���'>yz�>�?ܝ>9Ϊ=?�?HA�=�&���)> c5��<�hS��r�f��?;�?zR��vf�a�r?��~=�Pm��'���H>��M?ma�>C�X�U�/?�� >�+� ���vG`��j�x'���Ҿ��>���>�v;�p:���>J�P>(n�<�������=��龒׽�'=?+�����aM1>!�>x.����E<o�>�?1.*=?��T������>GC�tX��P���+���n(�^i�XqO�Ȕ޽_����8��������Z�����B�>��,�$h(?������=㨆�|8�v]>+�A���<˫�=�3���Mo�U0I>�~�>�rN>J(�
��k��>"���Q�����>C���
A��>N���l?��?k�=��Ӿ���>X$.>�mi��jL��o��d���+=�%?��}�!���T>"�>{�a���Ἳ�[>]�?m��
�X�$��e�;>��G����<�V=?�B?(c=�e���$D�=���x��z��#It>`��>LL�=<���n���q�'?��i���9��O˾a�+����>�Hþk�R�-���Q��f�c�>�˖�3A>|��>��?��>1�>F	��M���E��>W m�Fމ����>�[c>㲿��
��kB�m� ?{���e��Aw=p��>�U�}�=G�*��E	?��>j�m����>�¾�Oþ�\�>�?J�><w?H6�=2_¾~?-��4�ڼv����?a3D�%Lf��ʁ>��?��B�b6�=a6b�Wd�?(�=={|��,�1�3?�D��	ӾԦ�w;�>e)ο!A �0;���u�>!����g����=�ޑ>�M���c0�E����c>�����D��.m��L��㑿������<l��>�A���5��B7T�[Q�>xYƾ	f���u�K��=�??�ӽ�'L�[��=�~�>���� �>��ݾ"�2?0p�;v��<HV��k�=Bm>�a%��u��ʾۆs>��s�-gK?�X�Ø��24�?TXc���E��a;��<D�A�U���pj������>w�3��$�lO��S��}?h?�d�>��>	 �?=�B>~Jb?Tx?��?��j>;-?��>n#{=��?�UG?7��>m� ����>�>�0�>D��<�-/?�&��
��?ۖ-?���I�b��h�jE-��8;E+�> �>V�Y?���? �2�?��?�y>?԰>2Cb�M�����>�nh? ��>]�G�TZ�=ѷ��3S?)|Ҿ�����$��RR�>�k����H�;�	��uɾ����_'?�x�H�=<S�|%,����>ٶ�?��=�8�?k��>�)=gH?k�W>J�=u#���>��2?��_>������>D	�����)��?��(��s��g�=��?`������>�3 ?��=ҧ+��~��;�;>`�	?0aҽ�.?���>�}��{z=�R��ܾ�jԾbួm���ھ�R�?/W>�- ?)/�>�/�����,�?�!�N�M�R��>b4?�������N��?����f"��x��v��>}hq>�?M���
�	�͵����|;j楿WȽ�у��������W����ɖ��D�#C4�̆���歾���>�㦾�>1l2�;�H�3
�>&��>�� �8e�K��߂H�F?=��6��x=���?BD˾��	�\tﾧ�T��4�>��+?� �W�?�%5�>"�S>�n>s�����>X��L�_�s3����}�pf�=pi��\���	.?Γq��U�?T�ƾܛ�=�fg�3�?��
�����=��)?yf����=�k>���>�?9T=h��?��s��b��|>���FL���/����͌��W� >d��5���*|�=�>C\���(	?ռ�>���ބ\���>�ï�b74�/\Q�K�"���?I&�>闆>�ë>��.?~�%�����E��?�)S>��C��%߾I?s��,=��?+3>�?Ϟ	?���U��>�M��z����:?����1�5�>��>�ӷ=׽�T?Tb����=ȤQ�$pڽ���=B7�>۱���������Ͽ�@=��a>�6�ো���i���%��<ξ��6��娾���X�5���;?���<�?`
4�F��=��ʾY9?�䓾�^�>���>Y�>Y귽��>��ƾߩX>[��"�>��9?�my��a?�%<�5��>#�>ڶI?��T�|�=�|˾F���Q�>�9�?�����=��>?��L�M�?
:���=�JH�4�?�@#��?���>��:?=���>=G��>b)?�N�>AW=$�<��$?N.�A)=T���;E?��!�0�>`h�>�/1�m��;GR\����i����k$�4^/�>HG��[�"b�>x���+Y��$��,>�Ɯ�0�l�ǽ��ʳ?��?�@&?ߏ�>n��>����Q��?��>��ȗm?��?����v?��C>m��>1�X>{�j?�}>� ?�F�>�`?�j���\?�g?'�[:�28?�?�J >(@?߹�?�o=��i=R;��*?;?˙�c�3��Z�� yH�ޡ
�h)?�j?L8=��v>�9#?��(?z���h=~8˾�~|>JP�>e�?����Jb?RnM?r���H8>k#�>}���=_�a>�=$�8��؞?��
�>��>~�Z?�gN>)ؓ��H?�$�?�[�q@?��V?��3?jG�=���>��-?u?X�F?R�����?�y�?���>�Ii������5·?�u����O=�D��Q">v=������ �N�.%�>�|D�F �I;�r	���o�1;>�6I�R.>0)���=yn�+.�?Χ�=��>�
���B��wG���>���>ӳ�^����˽�:����(?���;7_M>�U�pKY>�:�>��-?�W����J��Ҋ>��(>W1��!&E��a�>�;�~�->�����r;S��=��p�ξ���H�� �=�;�Y�W�+='� ?��>�+ξ̬�QTP�m0�?,���ք=�nE>�>��V�Cd?�(ž���>�sn?>r�>a�׽&�Ծ��пM����,��ȃ�>�\׼�I=�^Y��h𽮆�>�c�=z�>�=�;�6Ͳ��/Q>�.������f㾔0�>�d�;1�������G@?o�K�#28?�1��SྋZ����x���f�.q�>:{)>ps?�u���&�?Dl�>��S�S�
����(�?P0L�7+��E��N��>U��ӷ=ꈽ��X���>���>ٝ����s�z��>ݾ���>�=������N+��� �U4�lO�����'8�����V=�����+?�\���xV>~�s��$'?ёr>�E������S-?<�=b�����>S^�>g�I��\�>��S�5��?Q�f�E��=����F�!?^���*�G����mC>w�?^A���(��cA�Y6!>f�r?�-˺聳>|���ȿS�E�/����>�!�58>��M���+޾�3�pt�^��>�p:��#�dV2?s_���qY�>�(����9�>�-����>��Ҽ	�~^>%O8?�.�>/�q����?��>r����̄��2?T�<>��=�Ȟ���1?�
�>�ܥ>P:��8�?��.?���>�1�>f�
?�ڵ�Cn�>ѥ���v�=�T�[��?��
�n�׾���>�i;?0[�>�R>�5׾�u�;��A����>�S��o=?�����/>������?v½�ʾ	�(��U��*?I�9�ڦӽ�=�>D|���{O?_��H�>E�];z�p��;둽=T	�����
?�-�>� ?a��=������$.?�)��aJ?�&?��|=�����i>��ý���> �U�g����?xʡ>@��=���=L?�d
������>����8���)�>���C��Q�>�6�w����-=���{y	>�b�?Z��J�y�O2�?��>n�8�;�r]m>Pn�>�Pj>��|�����i&�<��?�70���=#r�+P$�WvB?(<?Õֽ��>�A�����+��>�D>��뼾��=ͣ�>֥��>��^?ĩ�Qg�>��>~KN?(��?	����>��$?�j[?G� �����Ѵ>d"?f�'?@��>0j�?f?���>��㙣�麛?����'ld<�+�=բR?�ܻ�镾y�t?��>�[? Bs���E����������;����~?���K?���|d˾�GQ��V>��!����EǾ�~۾���>�����}D��(׾�8����y��g3��И���>5�>[��%z5����:?��
��[ӾE��C����輠�*=G��>r~���iM?�0��@�?�,��Y�C?K,�$WǾf�+?ҹW?f�T����=��?�_�=�W�@9�&��h7�>���<p�$�u��=1�>Z�o>�&��?�Q����>H5�^_�NY>���)?�Vr���"�����?�\L���I&��痽�~�������<��i���sʿH��lɾ��>��7��+Ϳ8?�[���˾��� ��=c%E�b�6�O-��?�8u�>I��{�D�L�a�>9�>m�<�ZH+?=�;�u�=ޞv=��>�.(�5���e=w�������O>Eh:�n��>���<q�RcL��f�>�±�P���/�h��O=����UB��O1�*5u>�����Z�N2�=<�>�T?a
��\�l�Y?nM*>�H��$:e?��Ƚy�b?p_�=�37�d(����>_�ؾ�wV>vKh?9��=�n���P��x�?��6?����>A���Vu�?,~ξ==�ڶ� .��.]�:^��оVb>q�/�_��W�>p4?�Z�{����;H�����TT�\x���˦�ps>� �.Cd��美�>B���kʑ=�B�=��>�L���*@����k��=bw����^ϑ="A�>�*m?�'y>v݉=<�L����>Ż<��t�I"j���>�p�=׍��U���񇾳����~G>4�߾/��W�O��<=�~?��2�P)��Z�>bC�=��(��.�������>#W��fݾ��;�4?T���T!�ڜ�>�4>�ޫ��\�	�sܽ�?�?��>�=�$
�>�)?S��>-�*?'r�>'h<?��>���<M��=��9�]�?%��>�m=>p�{=���>q_�>�S��pZ>���>2�s�/�!��澑8���ѧ��9߾W (?OGU=�t��u�D?�*�=�V��߮�, 5��Rh>��D�p�h��C����>��P��9ӾC�=�cD���a>���>��>�
$��E�������?�s���$=JM�v'�<\aF���= �>��v���!?!3?�(ݽ�S?�^��QQQ>6�@>�A�>Hˁ>=}�=�7|�P���G�>ak>h�۾ %�����a�>��?_�^��!�<��>i> �%���Ҽh�?F�;>2:̾�E�{᯾Q����ھ7��>����n�.�O��8?-� �����콻��>,����ٴ��^=�AM?i� >1>��>N/?�Ҽ�ϖ����i�=�QP�7x��7�7�׽�>������F����=�]?ՍW��=�U�>�ξ�/�� T>�t�}�>��&ܻ8��>��d��F�={�I=�/J>��żZ7��!Y����<��a>�p?kS��0���+	=˻�>����@�̾�=k�i ?�s��3���(���Ȑ?2K��y袾NW�>F�1� O >�p�>h5G����>{�>Gn'�t#���M�>Yr|>�L�_J���g�Z�&
��q
���?�BC�����.Q?��^>�t��ԡ�^T�>�@�>��|�����0� �&�>�5oz�#=k>.�:?�}>&TO���?c7��ؾs��>�A���qI�O�m��{��Ⱦ�f>�n���Z������k?a�r�����?�ƽ�������.�J>M� >��Ⱦ�_��Xs�>��>�{�<t9>���>�`��+�!>��<.�,��@�>�5���`��ѷ�>�xI>:r����]�B>��;i>Ͻ�":=���=�j����>�� =��=�⼀I�>�˽���>�f��I����>�5%=�g<���>|�.��Ԃ��ֿ?���&��>C�3�z�ݾ�؍=�±�4	?\��: ��'>�Ǝ>���� �ݾ��?��>���>�X��s~<>��t$�>��g�>�~M���|>f5��a�>�����ޓ=S�y��ON��}罨��*Jn>&�����>��޾�˽����� ?	\���q��`��s�>B�<�?��B����:K����g1>�M�X��=��b>��?�W=���=U�=�D�>�9��|��@�<3 �=i@��$2��m�>���>�N�[�o=�V�>��9>����7T�<�H�>Ќ��ʦ���牾�V)>F$�=�o�/��>i���Œ����>'c ����������mf>z�,=i�;랾!}�>��>���>��>I��>>j)��݀����!�TU?�4?�,F�b>ڢ=�><� >+�b>,�?q��>2��;�F%>�V���1	?瀀?�3g�b&ྛ)z>
$^>Q�`>XѾ0��>�C?>�����t>hN�>��Ҿ]`\�ͫ3��w�<�|˾?G"?Օ?�ᘾ\��>�]�J�=��?�>�۽�2�$�0=����I���>��N?�J�& ��02e>���X��>v���||>���߾o_� S^��jb�4�>����㫾��?H+@?�H��G���yV?��>�/��&1��kŀ>ۭ>�I�=���p�>�C�>YT�py?�*J�A�1����>G��>#��IU �Z�>1�>n��bIv��ֽk�>6l�Zr���<�>$պ Ỿ�z�>�rq�2x>?��==�,>c�ٟ&?K)�=rh!�&e��� �X@� �c=F���I��s����=Y�g����=�9C>�/>�e���$��iZ>`�?�.�>�������=���>Cߗ=RF?���=��r>�<?�6��b��7�Q��>�I��ќY�2����>�&�>�+<��ɾ�%>��?��!Q��I��nھ-��>E�ݽ1�p��8۾�>��u>>>s>��9�J�g������>�ܫ>6�9��d��U�>�Q��F��P�={��?�ӾZ)�@z>��=��?��*��䎾�w�>࠱>wPg?à*?[��_��>�߾%��)��>61o���&�$���*3��bs���m?��?������x�?��� '\=�轋6�>.鳾c��=�K��QR?6������X˼K?�ξ��n�I>�?��M�>��>�`�)�
>:�'Rὴ.*����>&��=�9q��)��ڵ �z���g��^�R.�>d١>�¼sR7?}qQ>I������	��>g��߻�=��#��J�>)�>��<=�����>ӏ&?�Ip���4���1?)�>^���������j>ɗ�><إ��ܾ ��R,�>��G� _�f�<D⑽L�>?�?X
>ח�/o>9�c>F'Z���k�T�7��g��֛�����H�oet����L���R���S�>�;T���I>�ߥ=����9��=bQ�>^⣽)�>����I*�}�K�x�-�
=�iG���~?��%?�R���T��ź>��>���>z��<O>���>i"5>AM%�e�>��>=�˾Έ۾x��=��P>�$����v=�h��Y^e���?r�>�A��x1�H9�<T!�����;>Y턾���>�;�>7��j'?��=+<���)�C��>�w&>=��>�+^
���>�>�A����>.�C?Z-�=s�Z���9>W2<􅼾�9=m��=��c>a���:����<�3�>���>��r>�c>�m{?��>���G��>����z=��?��߼�о�Ǻ=_�>�a���yN?|p?�W*�gچ��=s�J�?����{�Ͼ2û�f�Q>o:��E�n>�za>��^���!���5�G�%�v�,��#���B����>��>Q�m>����=%�
>�.?�?[��.p=��S>��>D�5�;��>*a�=(����� �W���>�Uq>6^?��1�=[P�>L M����=�>���<X����J����νL��\��Eߔ�Rի?Ӭ ?գ��L��!U?Ѽ?�Y>��փ��>XC>nVP=<ھ���>��>���I~����J�:&?�s������?��>5V[�Kዾ#��8 �>Z$��l���E{���6�=�袾Zk�>�t����'��z�>:^>O^���̾&���Bz�>s����R�U�˽�9�>�B���a�_>j�d��k��a�>�C1�	�,�3�=܁�#{-�
ؼ�@�0Z>�:?��B�=��H��>�n>
�m������>׽x��a<��>��>�D���V����E0�>��$>R�������՚>�R+�����@�>��?���e�˯L?|��=�^�=�	$���?�7?;&o�kȾ2�)>�~ν�^��&�>䞪���/��W�>C:�>��
����'�<;��>���9�rQ�Ǭ�>^� �����G>^)?�����{��>�͞>�����e�W�׽��>���_���쒾{�?�C����	�>�2�I�>�� �>�>+H[���<@�t9?���9�ɽ���<P;0=w W>WUJ?Ϗ��􄣾m_?�eI������>5A�>�TM�h-�����dU�>���������$>_��>���D�W\g>���>��=�gN�G�A?��)���v�Om�>����F�>d�->�l$>��-��>I}E>S�ʾ�hԽ�W?���s�e�a>�>}3��zG�Iξ�iF?Oϥ>��{���&���=��w�
�8����>|:=?���ժU���>��#>B�����x�����O?Bhz��#	��Y���?c'�B��<(�>~;,�>�v���M�T'Ⱦ�G?�kǼ���Lwؽr_�>�M�>* >�#~��vW>��!���>f�s>�� ?��a?�z��Z�>� ���<�(+>� U=�gʾ*����ir>fV��\����=�-�<��1�cD�?˨���j>؋T? �>p8>��̻�W(>9�?=�=��6<m�d����=;�����$��㸽�3�'3$��O?5��>�6�>�@Ͼ��>�>��>��>1!�mR�>~f�>X�=9�=iʡ>W����IV��-?�#�)�i����>�	?{��=��?��?�a
?@@��i��{~�m�/�f�_5?�Ti>0n;�::_?xK<�qǾ���<�n�>���>I+>�Ǧ�L��>�g�=�fh�]"�߰�>��>�wR?��=qgv>��zB޽1
=��>���L�>�`H����=/B�q�B�GJ�>��0�s2? ��>5U>�˚?[?@��̯=���=���>f�n=��>_z���!?:=yR�����6c`�� �� =AX�>���:��Z�%?���>�D��P�>�?��>�2ܾ�
	���@���O>��6P6?�A&>,���R�n��ǼlJ"��ž�3�Y�\>w���_���>zn?��+>��l�?�#A?���2��,)����>�����o=������p?XK����r�<,�T�g?�_����A�x��>#)�� �c�>���mo����?xҊ������2��¾8�D?��E��&R�X-=��=�e@�76�?�A
��^1�2A�>�U�����B�}�6=�vӽ���`wF>V[i��o�?�(��$-�A6�;�+^�L?���9$?D��=��˾��>#�#�Z�"?< �>�^n?t)�<�EӾ\���S���y+о�9ξ2w?_���M�T��Ѕ?�1>P\���*�É�=,�=�C��A��d�.>�k�>V�%���N���>b�k>
@� �>\�|?�վeu̼zt��ֆ�Q�>��_�
b�b�?0�>�iԾH1���/3���>����j����>m��>���Sjؽ�o7>��8��;��DL��b >��V?��=!���ᖜ>��?j�}?���A��>�tr��٦�9_�?�X�=&��?e��=<{��y���w��p�>v�=�@?�J��OO.��b�>Vq�>��ʾ%pT��m�=�_�<�꾡�I?!e>7�>ş��}�>m0޾%��>�Q�=_?{�+�I�D�Q9>�q�)���?�}�*�<i|�>I���Ӿ�1�=)鑾�7?�����G���i?�����n,>׶�>uz��.4�M,=X�X��1?rA|�R
*�s&���8ͽN���m�?�!�9F�Z�ݘ>%�?��۾h��=uw�=���gD9F��i?$҉?�G?>E�=?>K"?��a�3�оWͯ��"��+�h��'?Ψ5?�ݔ�̫��d�@?��>^μz�����k>&Db��oC���Z�aD?9!n��JO�َ>�#��[��>�=(�>�a�<އ[�7!�R(�>؞�����w&�>�^���0�P>d?�l_�-2��zT�>����2Kw�� ���&>�->?^x�>��D>_�>�����9sw��y߾�6�> nR=t^N�U��2�ע�>� ?v1~����>���>z��>���>�{���U�?�v>P���#�c|>�f>�R>d@���>��); �оp�ǿ��>�<?e<:���f+>JY�=����uK?�z)��3
�i׼Wm�ߕ������=�*Ҿ��>px��/:?qX�>���>�~�>K��k޽�q�=[�羦Hh?g��>ȝ"?!�?�S��������q���O>_9"�ig�?�Q>�h�颧�e�>��\?u?5Iv��E?��¼@�>`OB��Ɯ?_�Z?�㶾��?�$g�U�޽�b ?���>i��� ���V��B����g����i�=5
?L�C�c���Y�>���UP�<W�>$)>��S9���?��>��,��
�>GT><v�>��9�Rɾ'S��ʢ<��p�ٻ�T<w�d��F�g�=3)���e>�D�}j��O���>`>O�����(>�J?})A>�̃���������P�>1.�>��!=�ND=Y7E����>����`[��ml(��K?���=oe?�>S�?>O���(>�7澫����fK?q��#��>[�w�/>�N>��>a5��d߹D��>~�>g�}>w�+z��w���w��T>LC�=� M�2��E�����i͑>�;��#>ZxI?�n�&�q�(3 >������>�ʾ�Ӿª�>���Z.6���B?Yr�>��>�Z>��z=�<����=z;�A?�䠾?Ⱦ�t���><-��u�>���׼�.�> qؾYA��Y}�IF?UjO�J�?QGK�E!Ѿ'�?��<-辟���=a?��U>��?Mz9?g�=(R�v+y��|澄����l��Z�>:���:�M?�>雽��j�-�����?T���
}r�I˾�q$�>o �>� �Ϯ����>-�W?�I� ��ʉ?!H>�,�-��<{�=�yv>q�;�@ž��>w
�>�S�������?�Q,?��佦1^>(�/?;7��&�^?�cg��A�>Gž?�=onQ?m��{D�?����T�!������>80�<���B��=�g$>;ϯ��>ܖ?_L?K�>�+\�L堾�tZ���ȼ��� ��_l8?�Lp>��;��'�܄Z�+&o=S��>Z�|�>�����>O����s�?nk�>=#�>��>�L�?jp����=�C ��վ�2w?V��>Wi�>��?+�Q�����z���ʫ�<�d�>Q��>w��>���!��c*?�Հ>ƍ]�P;z=[�?�k�r�+�T�2��!K>a��>Y���o��]�>��G>]�~= L�qH�>�s�>ZN��������=��= m���l2��pl>D�>L\�>��>�:[>�����n�ÿ>?�Ƴ>��G�^k?H;����4l�=��q���>T�R?� >*=�F���(O��ý��?��>��h��<�����>�T/����=/$�>���>
d�>�Ϙ� ����w�7�J���[�"��;�1?��
?"�w>��ཕ˓�/�i=lM8?���ւ>$�׾�N�>�߀�{�=�e�>t����ޯ>��E?A)�=��>����*?��)?��O�e!>?��-?Y�?�X���,�`���9��l�7�]�����?s�=�������Ҧ�>�l|?e"�>�	���>���=�eE>�����?#�?1Ğ�xZ ���=T�
?�_�˰&�@�V?BX+��ξU�=�L�>:��>�ᙾ�S�4�>|�=�y���@?-O�W���^?���>��)��,r�*��>��>��=�Z��=�?k+���h��I�>T�)��6g>��f�HIf�_L�>z�>�َ=#w}>h����wX�>QpH�1	����??�=3,.�S��W��>G;���E�n6>yio>j!�>�녿�j$��Ub>��>3sѾ���d8?r��>�0C�:�;��`��\���A�$??�پ4R?ZS8>^֋>��	��,�?R�����0��!��0�>/�>�����X�>���z� =fd�>���>��@�]�e��py�>�H��]λ�s�=���>�	����P��L?]q�?��T��~��!?���=
��=>߸�%ё�Ѣ�>��!��t-�:$����F?�M����K���f=��>�b>�)���?�	<=U�_�'?�s�w�a�;��=���c�?&��>]]�>]��>ͣ^?V,�>�SE�[S>���;��?�󪾖2����h�g<�ʒ��<� ��c8?]y������'qX>�?�z?箦>�󈾈��� �3��;Q�iq���>�c2�>q�>�, ��ﶾ45��-*>�@H�[�e>�&�>��P?+�>�$��xe���>]�X�>&�Z�ꆫ>�u���w�J����?#9g>�5Y��ѥ>�K>.~=�B��u���>=>
=��W�?K���j�?̣��@��MR��/X���R�>����`?�R��E�>�£�i��=�� >�ټ�TH�.�����_<N�j����� �O���;R>=.�	?��^�&
�!N^?�?�>-!�֌�>>���=�?�Q��2@>r ��:{O���a>%�����u9?��>W��`�=��e>z�?S	�h~�>������H>k��*(��󉊿�,�>�l?b�'�d�>��A?c�.?G�J��_?��>V[>F���ĹV? �f>�>��C֍>;��^:�>b���>���=�mU�ȥ�=ZB�>�	Q���>G�]?��?��2>l�1��dm�ؿ����0��Y>��>�G����?�X	>�Cs�����>;�=L��E�>r��d\+?�e.��9��4� `@�,�?�>2�0?��^����<�=���^8?�*���>n�>^�>�@¾�&�B����S=�bc>Ո�?�>���?D�޽���=����?>s�݀_>3�Ƚf:�>���>���C�����+������⸾7�?� ܾ�9���wz>���>��꾷ă>�$F?��+?���>3�����P翾���<?�꽾IX��Qt>���>h$��e</�D�]='�,>�Q�Nr>��m�[� ?��>��>pK���>���6�4����=Qu�=̴�[�3��.���D��ն$��#�<���>:ʮ>V������1[g�tms��7ƾ��`���ɾ�=�k?�>�.}�J�}=�>���$?��4��j��P�>���r=�����>�F��:���k�>�>)�Ҿ���K�(L.��؅�����:�%�T?�GQ���/���N��%���>=��>�W��m������>�j=�����>M�>�{?��>,m��g�]�1vw��#��z��>50�<_����?:��>������,?Sm�=�f�9�q��Ø>�K�>r�.��蜾�V�a�>2Q�>\ ��YƩ?�=�{x)�ޙ�>�N)?�h=���f��Z�}�0��>(��=L���vԾ�f{=">��߾XJ?����ɀ����9�c_6?a�w�v��� �p?�Z5@?�L?���<���>��i������> ��>�7�>��%�U˛���S>`�=f_4>-c�s�7�
�۽�I��g�:﫻+�F����>O}?��@9���6?t5v=Z�=l���Q�>�ϸ<߯r?d$�����������>�w�M����	?�MJ�|�;>L�>���@�=׸����>�gd�d«=�lӾ*z/�q���43`>���>-O�eR�>_q�U��>�{�>v��>2�q���>Ir?5�>��_�F���>\�����+>��?���F?�m�w��=W���|�(?Y����阾
�¾�ސ>���>�==�sE>�aE?��?oO
���R�i�tƩ=�zI=�S?N��>@����?k?K붾ә � M>�/N;��9�_���Y�����>�4��/���F>��>�QK�R�>.��>Ci�>1_�=ۚ��6+#�*�>?f�,'4� �>�N�J)?��>`ν�����L�>�f����"N���;��?�?��>���>����)o�=A�ƾ�U��8�5?K�?c����2>]�=��h>�=V�:?p�;�C>hb?i��>��C��I�?�X�?O�̾=;i��?���>��>����~F<�.>&&>?�mh��-?=FI?�ʗ?�)��hO���=�zѪ>m�O?оj�:�0h�>�\!>��M�T\�>.?�� ?�?
T�=M�8�w��r5?w�?���9g��='��s��>��>Y2�><�l�ұ>;�}F��+���@T����&wG?��g?rC��(����>]��> �!>Cq��OqU>�]�3��>E[���Z7?�d?�<?��<>n���΁��	u?"��>���<*4�Y�0>���=:{A���սL�¼
z�>؁��ܾ����~�a=+P��{�	?�	��s�;�\>1�??Pp0��e?2!�?��?:�1>�:��V���+�G�f�/{ ���4��}�=ɘο�v9�H�>@�>�O��|J�%q�;Rع������B��J*�>z?e��>���>�=�>(�;���o>i���"�c>�#���=��Q��J���z9���� x�=jx�����>��X?�����u�&2������MoI?�>z�i��������>�\>D?�ꖾ��-����>jX�>��=]�����2�ӛ�=-=����=�0m>�?
��1ؽ|3=��3���D��
Ӿ�?�Q�>�KO>B�>"�?�Mt>;�^>[�ɾ��Ծ��/ڗ��s�����U�a�Ƚ"mW����)��梽5L\?�a�:�����>���>\i"�͒�����M��=�о�ɘ=w�3���E?�r�=��9=����gU�����jd�> :r�l�J>Y2Ҿ���­ν7`,>��d>2���4>}/��U�*�$� ��h��H�~>u�$?�O��!�O?|<:���>m�B��[x?f��=|3%��2B�@	�>J:�>�H��3����+>C�>7Y'>��S�?Us>�8=!����h�>���=a��J����x�=��-?'׆�����H���X�>�Ǥ=�,<>> �>A�F�8?E�S�>+!?�=�F>�X�>�®>�w��/����⾤%羕���0Ծ��F?F;�YRB>|)�>�3>�V��ȉ�>��?��>�ĳ��c���J)���n�M���M*��q�?,��?�=ž�F���Q+?�>g>��>��_�>���=[ ?Dc��@��>�?�o�?=�龠����x�=C��<�?��kL�W�>i��r�>���=!{>�P���#A�T�!�R�O��,���!?e�u�7�d?�(>�[>�jS��WZ?&u�<6XV�ў`��R&=��>hyk���n<�>y{���?0�%�	Q�>1f?k)��{����?:w���1�WQ^���ӫ+?���>�,?7��>Ok�>X��> h�=i[G>7M,�?� �҂�3
���d>?��9�>��x�>r8��#>�<�v'>��L�����>pٶ���N��*��B�>-�����>G�?k�?k��=r���=�=M=��gq����Ɓ?��2? Ro>�G���[<*����;7?�	����=uT�>��H?�˄�π	��y��¡>���=�����~н� l�A�޽v�D�x��>�(�>O,3=ET?�<�?#	�>:����r��>��=�|�վ�?'��?A�L�Bݡ�*�;H��>�Z;=���z�>9��=fث>�@����9?�L?��J?!�	���ྭ,?Eq����T�$��� ?�:�y�=<r	?�i�>רt�ԛ���Z>�5H>%hӼĕ�>/N@�`����^?ڮ�>��%bX���>c0B>Sq����ν5f���!?t6j��j��k���P��S?n�k��>���n]C��V�x}��TJ2� �ܽ��>�q�|,���^�T �>�?�V�>�%�������>k�ܿl��=�9e�YrJ?�3��^z���|>�7>X�{�����`�v?�#�>ߖ�>X����o?y�>�~n��+��!,>1*�>�=��V�<�&?�������>��\���o�½�%8>�<�>�]C��q���F?�:>/�=�Ӿ1�H�e��>˂��I˝�P���c�> M�&�j�|	?���>���՛q�`�L?�,�=|��a= �'F >�$m>�j�j��>�l���	�>o����$�iE�����O�O?a,�;��>�>����K��?6"?�~�p�V��汾��e=���>��>ҿ>%G?��>z1�x?��V�>c�>W��\��E+>i�>��*���쾎�Ǿ6�?��=O"½� �Jj?��r>�s���d?�����Ѿ	:?"��>/3+>)��`�>�ku��a&?v�>�i��B�r����>�_�r�߾��>��>ީ�B�>n��8$?01���1�=>T��?� ��;K��7��<p�>�R��ο���>RҰ>k0A�G��'�=�C�u�����|�Z���*�XF?�'H��L�sB��QBݽ���Ͼ��d�	�c}�>=��=��ž��`�hh_>�?;tU�>"
�>�O?�N���l>��L�>����<�?ڽ?���=����)�=��>͏��D�K�|>��þ�</�d����Ҿ�AQ��2U?%�H?f>Û�ZS����I?�C����>�n�>Nf+?Efq�ql&����>�rn>����½Uz���Ϯ=)�ؽ%E�>�:>diS?LV>J$?�ϴ>aQ?�� ?
T$>�J=��&?�jl>�5L>���=/B�=lI�>
���SŽ��~>#�c?�n?1�6>ԟ�=�~�>A�5?{�?y����Ծ7!���z���?�v˾VG��b+��~�p?�[�r�\�KT�>#�>��F����Q�>A֡>Ǖ�;6:���A>�i.�u5����澑�)��q-�I�>��>7����>�����q��1���a��'�p�9b�?h?��>�=�>�ֈ>w#�>���\M=���=C��>v�>�쏽�?��>r9�Jjr����>���v��>�|����2�\I�����?�>|�>`�I�t�?�m?<<���o>��wI�%�'<7�`���E=o��J��>�>��}#?�Y��AI�3>J�>&���?!��.Y=.�i>:����@>Ȉ?:;�>4Խ�h�Q>��	�b{�?P�v��pV�(_���>^1Y��`���w��u>`.��h(?^� ������f>a�Ծ�B�עѾ0��>���u�	$�Mn>�$h>��¾�H���J�U��=Ve� ��>�ʎ=��R>^|$��ْ>�b1�&݄���>�xr?�L��d��۾{թ? �)�v\�>:�>������>�w'���/=�g<��4?5�E>ؤ�r��>h��?d?sW�:
�4Ց��2��,��� �>�)!�E�߽��ߧd>�}��-`��Z�>��? �$�	\���"�>��>��F���R�p��>�ڙ>��E=Ӝ�>d��=e��5�	��E������S9>gq>��>d�"?��e�(^��Ƅ����B�>V��U��>'V�>S_�>�ve�_��}e>�1���Y�����ƕ��D�>$$>���>/j�?^q��M�+?f�d�W.B�ق�>����a5?�?��)?���6���a7�Z.?���2�c>6��?nh���S�>p���A>d��h?�?4=?,��7�Y>�ܼ�A�=�hB��̼)�6��s��)#Ⱦ9��� ���Gܾ���?����t��?�c��o��Jվ ��O��ty�n�I��݉>f����>���=�o��#,�Q;	?�sZ��up���=�D>N�n?�7��
A���>L9?��"$�>.�Ⱦ�'�>��>m����ބ�'����>�E>!�_�`7��[�>�-I?;��>,��r��?l��4!�>N��-���o�轃�V?�<{�;�A���[?�`�><E=�=��r�>�W�>}��h
�M�?1:���>og��Hz?Z��=�qh�����X ?n00?KJA��&��+�,�؏%�V�>�j ?������>�	8>��>X����ϾNQ�>�� �����y���X����>V��>5d�>���?`!y=�j������h�<�=�>4K?4�>Ư���<�.1>h�>�]�Qn?��~>�z�=H��>p���O�.G�=HQz>k�/>C�>�`�>|9;���G�t|L?�?�(H�.�h9�>�8�Hb��Nu����</��<C�2�s����C�p?I5?d-����;�Ƃ>>ta���4>NzH>kξ��h=b"�=	�(?�ꔾ�푿���c#�=i�Q?��>s�>B�>��>,��Dn�<�@�>4��>Z� �̡��Zj>��|>��߽�2=��!�?���>6@�U�t�*��?{%?���c/{��d?��!�Ë�>���>O��������"�>S����߾>a�>�{�>G���M�]��[%�=D�>��E�#ܬ=F�=�>	�࡜>���Ql;�5>0%>��d>T�E>��>�B�>�q?���Y�I����*\�=�D��3��嬽{.Q��ɀ����"�_><B9;*�L���徖뀽���<� %�Ӫ����j>���>d��l�>���9�;=���>�p�>���=���<��lQ�>�e�=�����>�I���z9Gne��[���/�=vs���P$�+�:���׽��">�`?�O�=m��<Z��8[��4����>	s����>���=sR�xY����Ob�Vp"�ן�>| >�G�#��R�=�Q�>И��ܷ�L��t�>G��6���F� �;�hZ��Ƿa��ӝ>>��;�i)���(<?��>�Ҁ��>�>=����^�>񺰿��?����wU?��>����?S�:����R�0�B�\?N�(�O�=�!���?-��;2��>����~=����/�h��}.�� r�v�5��;>��$�gƾ�i��s�>:����5m�4q�v�>,�о� ?��G��!y>^?�N? j.�!����>�!`>�����G��v׹>�~>�.�?���>F��>����ݵ���f� �?uɅ������r�>15?Aw(�v�����>�?�t�� �=�?Ϣ�>�E?>(�>t�����:?"&?�'U�w��=��J��>��?�:>�{Ҿ�v��?�E��J�>�� ��1����w>�ż>6;�=:�?�2>K> ��?qU��te�1J��Mλ�g�?���O���>Lя���>��T�M�?���>��?�$7�]&�>��?bW�����I�>��#�n��>�M5�x��<�|5�>-b�1O?�]�EN`>�9?M��>
����*վB���}�5>��>�=w�?.�?h�$���>��?�>�Y�Ѻ����`>�5�>�;�M�C����>�J�>螾\�Ͻ���>?Ѝ>�6� �>^	>7�=�B��
�U���(�ni�=s�"��D���� �P?xE#?��(?��,?�>-P�>��/? ��?Cj�_ʾ�殾����꘾"[?(��>@���<�-D=��=8	C��Z���b>rgվy��M_�Vة>HhS��->�1����=��#?C�о�'�>He�[��>sv�E���{>پk�m��Ӏ��⨽{��>�R8>2^��TM�>��\=蔃����ե�ׇ��R�?M�*�+�]?���Ji�v����Y?�_T?♬��팽{&?���>S}?�H���S;���Z>�1�hr�=y�?e�>��f�����[�?T��=�á�����퉄?,�>����O=|V'?�%=Ĕ�>��#��[?1��,���X�Zr�>�8"?�g��]�޾�,>�A?'+<6���!FO?ٹ�>I�d{�>���?����������>������f=��?�Z�>�`�������?=*�>T��tJ�;�}c�����W�_�1Զ�i���]�U����>g1�=�ü}~#�����y�6j�T8��F�ӏ>cf=���Y?�Ep��μ�>���3�>�3�>���딾��b>Z�>2�¾�+����>ʥ?����%R��k�&?�%�XV@?�5x�Bn?�{?���>E�˩���,?~�>?�����޾��y�RRL>��=�6˾�"��2�T>�+�>`wjm�^? >��??�{�����D>˘�>W� ����<�w�6�
?5��>�`��ZK�4�>��[�=1d�>i�#?�0��D?���B> ?B�'��=�����E�=}����<2��vC?��c�c�R���ͽc���A/�N^�!1>�;�=cgq�%W)��8�?���>Dv��{��=�����=�\��s6�w�ؽv~=��|�d����T��թ>��*�˼�]�>��?uU��O�>�qr>��?s8>��؎=��>�J>2�>?�.!>�����ƽ�bR��(�>��d>�]��_վ\��?8�
�7��b�����>2���~6�>$ds>\Il��Ҏ��3�9!񾃢j?�M�<��=�_S���=��ܾ��=�q侻�5?��I��l��R���9?:໾;v�߉����H�ľV봾; ?��1?�n"���Q���E?��%>l
�������,?�%>?��<��Ѿx=H���?�>'%��,?.�L�RG�a�'��>�eM�@zz>h狾(o>:r��G�5��B��I�>$$>������>��8�\5a=�1�>�{�K�¼�?�?R�=��<�����ӓ>���"p뾐�JT�����qn?��>���>���>(w!>)�J�S�Z=���>0h�>�E?m$?~&�>B�><.I����ր�=�� ?�C>��>��?d�>c�">�,$>Ε�>�5�>0BP��B
�� Ծ�.�l��b��<~\,����> q>�g�̐�=�����Xf>\�?S�l���t��IN<��x>T�����Y�p9��ף���ܾk2=���>�<=�Ⱥ��̾���;�Kǩ�[��˒�>f�)�	�l��<E�N9>�=�&g��@�>UV�>�����>�#>�T�>6�>໶�{&>�'>_�<��^j��_T��f�W��=��2<�ۆ=3��>��X>�U>I1%��z���>��S>�u��yC�X%ξ��|���m�?;E�/�������>߃=���d������>9IW<^��=�՝����>��<+7�9�K��z�>���=��$���
��������E3������>$�վ��ξ������>�?���G��� x�i^4��t�>��d��$M�˓,��'��a�
����>�˽��x��H>1`�e�?�r嬽ʙ����^�S?��d�w�J�=���1�>�#�;Hni�˪7�7r?;K�y�����i���\?����0ak��[�t���%�=�S�>Ob>���>~Y�>� ���I��X#ۼ�6?���>�*7�Â�������
�n�
�k�=��ʾf.>�b>_@=��l�ԛ���>�
�>eJھ똶���}>"��>·��M+�=bIJ=!T1>�伽I�=��>ė��scH>B�ʽ�e�>mr=��ľZT�=j9��0�x;���Iq۽���!�>I��=�� �ϗ.����n݄������>�a2>�6��k��zي>X�>��>�>���>G?�2�E�q�V�at�>=�/?U�>��ܽ3P��P�>�6�>�'��p���0����ht(>��G���A���=��ʡ>�T�>?���X	>2����Q�=>�ѽ�<i>ŗH>!O�>]��Y����fw=U�>-�<�s䎾���� �=��>[�:�����	��[|�����iM[�B��>�����[Mܽ���>eD<���>��=<�&���>�>)��>�C��\��>���>t� >�U��r>�(&>|�G_c��3� 矽0�����=�$�x�о�-ݽw}w>�+-�wh۾�x���t>��2��=*_"?R8>/ �{��>���n�ޱ>9�%>Y�=��=4�ܼD��=E�>���J ν�_�>#�_������o����>���>���<��7>/H�>u-3>����h>�r?o�U>8�r������C>i�=l~<u`�>;�9y��Y���5��`��)���|�>6��<(O �Gʘ�x�>���>m�=>���>�;�>}ؽ8l>��J�\��GŐ>$oI>�:>�&���^>�C�>̟�>��>>6�>fn�>�ۭ>���ת�DBE>�H�>�G?O���C2�����>A�>.�<�j >9��=��>Ֆ�Fq�=��>x�>�ma�j�>]��N�7��>����4����K2���<=՝�	��>�L6?���>ҶH>n=]�C��o���>kf�>I¤>(7��B���|��\̓����=��\��#H>%Gi��]d�[4�h�D>Zѽ���>g�.=�͗>;/;��r�����>���<Σ���>�`+>��=�Ÿ���>��>�F�=�A>BR��ȨO=����d>@��97��a�=q�L><Y��`*�8Q>���>X%��y��T=tr�<��	>|[=>��*��V�>ׅ�=�f�������>���>�l��PW�r{�����Q��h����w>�o��a径�i�\)��C�y�;�����h�VT#����xT����>�{)>��>�a?��?�F%>��[>8Ä�RR��>���>8�(�X7|��R�� �>�j�>OE�>O�>0�>5������������L�S2�>�F6��4�=�U־��urr>ɠi=��=c؂>�½>D����<���e��>��Ⱦ��辀�S=I 5�U&��M�S����GV� Jo��N�Z�:���;>��@;	{�=�b�>��=z,=!�
=�魾�m�� B<Z�?�?e�j=4��>���^��'[�{��<t�:S?��'>�k��z���œ<�NR;��>Ew�=�h�>�4Ž%җ��ξ��?�
�>c7.��!l��\�;ס�2�sd�>}�?]ly�����]�^���=�#>�>�=�m���O��i���c�ȱq����>�?y>HJe>�a�>��[���8�콴t�>1��ɢ�����X�>P�	?|�J�=[�>��,<���n4�>d:>�n~=
٪=�)�;�t=�8�>I�w��K��JP >d�^>!���������׃վ�S�Ѻ�>K_>"���G�<o��K��>�C���,�V�>�� ���p�,඾�&�#��=�x�· <Z�>>�����>]ZB>˧�>���j�ͼ�ꊾtXC=�*H<�P'��U>�,k��?.��]#>cS�>�5T>�����=���=�[>�Ḿ�#>�K�=�?�׾t��=��>D��>�t3�թ�=���ڪ�>S?�T0��5�?0侓�ֽ���>6#>R�g>�!Q�k�9��*׽��(�>��4>>A>��>�S��E�a�u���7j>��:alw��qʾb^>���>I����>�� >��:>�n;>�\��c@=T�Z	��m*:��<2D�>0S���Jﾾ{2�!�<	��>�Q? �N>���>⽠��=���B����>3zE<?�S�>���=;�>�^��y�`>N�J>�x�ϯ澘)g�y��>SY<�E�=���=S��=!%=ڀp>��#>7�[��=%žR��N������$;=��̓��<�>a>�>���2�O�Jtt��n�=�����7�:�<�B�>��.��^i�z�j�Fχ>�������>{��<7���zt�>M�	����=��>���>�?���@�XB`�ڏݾ5�7�����o�>���;ao{>w�V��:^�b>kf�=�s��ݝ�>��4>�=���4��>?"�>>�=�E���<��o��)ý��=�j/�- �>7�����о"0�>�ka>PQ}��BžER�==��������9>f��vX�=}�қW>��=N���.�a��>�X���2�����>o)�������u�mC��`��>�x����`����4]y��a�=F[þ�f,�b��=t�Cq络����<�y=�Ș> >��R��=h�F����&�k��G˼[�>������O�>	(��^j��	o���>y��M����|�p�N>��?��>��<,�>�YG>��(>�j��LX?�OA>���>�����n>B>���=ԭ*=�����$׼������/>�N=0[��_�r�#]v>����v��u�վ>���'�D�����=����=N�ȽX7>���=!TC�궼J(I?�����D=�qQ����>������N��Ͼ$/�Olܾ��<ln�>�ؾ�r��;ä�|ޜ<��1��t�J��>M�>�;�7���>A���L��>;m��<=�7�)��*>�$�����޼��k>h��2ȏ��O���n�>�\_�7�*��=$?�%= 2�>��ʆ�dS�>��Z��#	?�?�;,�α<�T��>�C >fh�3~����>9��<ԫ(��-��Q>4W�<㒙;SJ�����>Q~�����%��"?2�｡)ݾ��C�~a�>:s�U�%�&H�� �>���q$~�҆H�}x�>ϙ(�M���~��>��̽��>������(���H�E���a���5?�O>���;����;���>뽺<fX>�U?��>�%=_l)�B�>}>�>�=?y��>�=��/�>�T�=ӟ�=�i=Q4K�s$������ꔾ%��<�m`>.���#�>�c>�<��Ƙ>� �?_B����=��J��`� �oVi��� 뾻���ʶ�*�>��>D�?v��?"߹?�Jھ;����j>8�?��`��X�>��>  H?cT�ϻn?<��>��>|��>�~�>���>O�>	��> �t�,��>'�H��.�>U�0?}��>���>����0��h3��h�;ѥU?����Y��>�@�>�)���3��=�1	�m)s<e%��uT#�~��;�9��k����?�#�}$�>T����m��";����>��>��K>�,�����e��>����ɾ1��>+>��S>�/y���?Ā >��?�U���r�>脳>�,R? 
�rӼ>KG>8�>Lk����/콌0?��>� k�w�>�1ɾ�.z=0��>p7�=����T=,�f?��*?����d��Iڑ��N�օ̾��ؽ��t���Ǿz�|�O�?��[봾T�=>�<�>+��Z�J�:�="��>�?�_�w?;U?�BZ��>�8p���U?��<�� �0P��K�>�'|��5 ����=\2O?07���紾p&���Y�>)P��˽�TM���y�b�W>𗎾��<0D?k��>�ń�wy��V�=>nS���ݽ��?��|����K;���>O]?^|(����뾣�H>"'Z�˽��:a���>��>�G<>��>�پ�q�>h�<I�?V�E�͚�>{[<����?�n���`?��2�=��Q�ń�>hl��P���V�}i�>nҾ=�Ģ?j:>@�B�L�_2��z<��M�S����ϾkP�>0�پ�t>H�Z>?�>x?�V.>
�b?E��>�����=v<^"��u4�FvG��X��o,P>J���9�����5�-l?���)ڽ���=�B�>mK$�a����9��@>=Q�=ԛ�H;W���V?BMq=�{?	է>KE�X�=j}��j�����w?���s� ?�\Y����>�K�W�߾F�� �<���=y_R>b??��������\?z-�=�뾃-\>�9?��>a���>mu?s�>t<I��58?���V���<�.���b���4���<n�%,��^,�=��u� /�=Yu��{�I{�=�q�>����;Y?B�C��L?)77>�D:�[�>��=�8L��y
?7���fޮ��?�=�f��%�h=��'�B�a���0	>�r�X�-�>DY>���>��>x�8<1���lV�ݼQ?d���g';?+g?ZR?���>I���$�>I��&<�>� h�ͱ?C�$�8�o>͛�?ྑ��>8n����U>?�>~���7#?�Q���?����+��1?.���+?a?Y;yk�>�>Yn������Ŷ�>3��dd!�E�6=byB�v3�>UþBI)<70S<N�_1�>��?���� ��MK���)?b�>�6?���>�뾐a�ڂf�/>�|D���?̱����M?Ci�;_�H>^4!?�C=�4�>ү�?���>��>�f�=}�>��c?����X�����?�e�=��?6|N�"�<>�S?���=��9��>����=���=Z?@N��eb? q��͓����+�>-��:��?�> �=�+_?����P]?�\�=W�վ�q�>{��ި<���bq����?�6�77'?�	>p`��ͮ>2ť>���<(#>zj'>v�b>AQ�(<:��e�>yQ�v=����?B#̽�ĵ?�,z���y?��?R�=��r�/E?6n?Q͌>��=r�92�=@ �>"�̼|j�|j<-�L���>.��"�K�S,~��>�c-�qRZ=T.�=
1>��>+_'=/��͏>cGe>�W�����5o�>,�>�??�:�Z��>U,�P&Y��*��r�=$����Mg�{Y��>^���3���L�<{�>&̟=�H:=W����a�>��>�>=Hw��1��`>j#H>T>�O��T�s֌�^?��!��}���X���@?��t�������>i&#?�%l��\���秾ۘf�e	q?�$a��I�>L퇿�s?*�y>�<�G��� �?K%#?�=ͳ�Ƀ�>�W����T>p
v����2��R�c��'
?B�Q�%�L�23��5�>P%_>m�9>�v(����=�����?;~���=>E��>�3�o�>��Z�B��>���>�*�c�O�9�����Ɉ����?59>���˖<��?�徽_�۾K�Z5?�qv=�Ǿy�W��q1?�.�L�h���6>�P��^]��N�]i��͘���?�Lھ��ݾ��
�s��	dֹܾǼP������U��gق��޵>�*?��T?�i?!/�1�=������9?����w7��Q>�@L>��ͽ>�X>�:[>�J ����>�:ʾ!q?B<�>jGP��1=�������h�����վ\� 8�@��Y� ?E�*��?�1��E�>�+ ���Z?2��	�=�"˾���>�ľ���=���	��>xX�z�>��!�
�}�K<D�f�^>>�D?���椟�?��>٭�>��Z>5�_��*��1����+��Ͼ��ݾͩ�l{�>/M=����\<?Q�:>�&?Rx����Y?d+?�f�>�ea�jO=?�S`>�̝>�����}J>k�����E��ڝ>Ǭ?�J?r ���l%��㾢=.���8>��F>X7�oR?_��>9�
>��>�ٺS_�?sp��A퇽c&�ݑ+=l_��፿�k;��ܽ�<v>H�:>�#~>�f$>�Ӆ���͆þ+s�>��Ծ��=}�W��F�>Ke�����:��Y ��� ?Md?s`�>�%?]h�?��=��7?��R?-������MД�ǫ�?(�!�L�?2�>�
&>J����l~۾��7>���n��y�	��+v�u%(�)nP?�j3��L�}�>�5�>�"�=S떿�߁=��8�#	Ҿ�Pe��q�I�O>K��>AK*>%žA�>���>�5�>�J��s+��0�>��|�OO�G��=<>]
-=�l�:��:?_�H��b�G�?��'�8��?��w�h�>;�|?�)�>C�T�&�a>W*[��C.>%�=����9�p�=k5`���վ���?t��=�i?z�G���?	�[?��>r���xY?f5!?Ǜ�>����~���HZ�G�u��Ѽ�s�>,{�><hK>�}/>���?��>#�L>_�����ջ�n��^?v�.}�>�Ų>ކ6��9�=��?=T����2>r���� k?3�&���F������H?1�2��t����ܻ}Fj��D������8�oq�]���9�ʻ=���!?�A����>z����>l�?�7B=#;)�>xX���M������k�yB�>�;;FF>������9?z&?ew=W+�����=�>��L>LA���{���>a">��a?(��Z,�y�
?��>D��h��>�r?{}>�R+�S����?H?n���?_��=�4ɽHJ={��>��ۿZ>D擿0$?tr���Z�	�p�s�>jA�,S;���?�k0�>���>�Q��̎>R}?��ƿ�=>����>����r��k*�UR:?��������ߌ�\L���j=�N���>�r�>p� ���>L%�P���� ���)�߉�?��9�Q�"?�-�=#Yw?}\�>�n7�C��`��Ӓ�U�����7(ᾊP?+
���������?u<���=�?�>�	�?�U�=)1 ?l�C?�D�>�9��[��>wM=3�=�0�>ko4���?���=ʗd�.�����%>�̚?�uH?U*���q�=��>A[��TLN�ȶ���)?%�>e��bS��x�=[O���2�e)1�QS����>�Z;�ſ>��b?�ű����>�ޓ�D�?�Q��]o�����aձ>Ӿ>�OT�J�4=&&?�p��N?%�\�:|뾧���꾾C]�=>��>�i!��
J��E�=\u,>4aT?�>K؃>e�T��%�>���S��>~r�=�oF�~|d�7G?����W�>MA(�v�=?M%\�\��=N�!�+��ځ>0&޾�1?�ӌ��}ؾ_qo>���������&?�n>�a��^���?���'�����¾Jy>�=ևF�ms?�ϊ>Ƅ
�m>���U��>�&>c|�>5",?=��>S��>+�>�}��k��[�?�?�b��*�g>X��> .�>L�?��?�D�>F�c��[����T��>Ǿ�c���*�>�"��"�>��>Nݠ� _��.\�Y>/Ѿ��>�]�>x�=p�M?�w>��S�6?�d߾"�r��U?<3i?�!��S��}��A?������=3��>�̳�MI=ʤ�x'?�\�>�������>0?�2�u��	=�Q(?�)�=dV�= �ɽx�����?�����&�?�T?�ܠ�[\�צ>�Xb>L/���������=9�v��=U|�>Y�	?\��=�.����Ƚߍ���	�?���V(�����y��?I�[�<�:�v* ���`>�I�=�P̾�Ҧ>^��>w?��1�x�j?�XT>�	�#���d]U?8]�� ,�x� ��??�P�%e��n.����>�a?Ծ�
�=�(��M�%>fت�R<ݽ2��>�¾��k>��ﾛtS��c���?k����Y������c x�g��>F�v��)�}3���>��^��>,��v���"�>D3r�&�A�j?�(�]����/>V���"
�=�n�=Ѣ9>��8�	0�I��G�l��5�;�>K ?�=XX�34>��a�{;�{'�>g$l��v�>�5?A����6��h��>f!����=�*S�2J>�fn?72=��(�.9Q?;ԽUaV����>�d?����#پ F+=
��>�Mr>�#��^L'�jZ�iD!?s���J��ד>��@?��̾Z(�����>%e6�		��Z�l>�/�>��ӽ�]����0��۞>̔�?�{?ț=(�L?��>u��'f>�d�����>k�ľ
�'��gC�����	?�\�=������P��(�<��Û��Aޥ�8�U��{?�Ѕ�	R�7,ž1U+?�M3��8%�K�>G�>
q_�!��@>�����XF�{��=h�<�y#?C��i4�������=�%���y��J~�3J;?�6��N>eL�>��>�.�B��>1���2�Cd1?�Z?���>�>I����>���>̀W>Y$M���}�W����>z%/�I�>�%���ѵ���>�5�n>���r����?�������j�]���i?�R>CA�>�I���$?]�>ȴ�=֋��a�-o>�fl?�Q��\�<��禾�i�>��?�s�N�Z�'��P��=�b ���P��*�?^=!��\x�a$\>]&�>l*�b����>�.`>�
�>i�R�:X����i���=A��� �;?�>��ľl�W>�\�>Ў� ᒾ1	�>z��\��m�0���0?j�?W�?�>�sA?� ���^=�A����B�)~�>�>���=�F�{����]�>d��=FTq��#����>bp>{�������?dY�>{�?�C%��xپE��>�*�?P��=ҔԽ[��>W��>��D�j��=M�>4ؽ����2�:��#�:?�3?Ҫ�>.����>��{���>}�>|J?-�>S�ʼ�+�>�2�<�� ���?�Ϯ>�?\�D=h�T��'�<��X=W$�>�ֺ=>M�=���>�:�v�=訁=ř�|bнW�n?�V�=R�=g.n�]���c6�?P�>�󲾶(:�4�6?lކ>y�>��P9>�8�>2X�E��=_�t������>?��=?ꀾ�XD��wQ�'4��*# >�꾋Nn���?e�[�� #��G?!?>�X�=�]>�1,�4A>>5�>��?��P�|z�>&v�>D}
?��+���۾�5� �����48�=$�>�J�[�����>��>�d	>� �v�����>V�P��P������
��>��M?4\:�ũ뾬~f>��k>cϑ=�ꪾ���&�>��d?�h��7r��.��[��>;}=�M� i�=,��>�?^�dO�������{��#?է=>��	��ݴ�~O�>�#>�.>:��=mC>��=�*>���*_�1�>g�����؏�>'?�5�>^-�]��Ԉ2�o�w��Y,>���e"�"�Y? �q�Y#=04?�4|=��J=q=�r��U֍>
]ž:X�>�f߾�^�=�� ����5R>w�\�Ѿ:�?���=���>77��"O�6��>t�? )����>���=��ʾ����%��>�=*o�=���=ewӾt�R���g�w���=L,��
�<]���<�u<eP�>���<j� �� d��.����㾌*�^��=�=#?��3>:Z?�*���3۾ �6=��>^p��̏r��?���#�>.,O?�D�,�i��?�>�䯿]�>m�> 鼾�f��N���gƽ萾��>3�>>�u߼ 8.?��8A(�\!?�K�I�!�ٺ�?=�?L�M�:d��B"?2g?�jY�N�����7>?@>>�g�u(%�5�=�5;G=�Q�=�i>��Q>I�]?�iu>|�<<i,�>�|཯(m��*=+%?*q�<z�v_���2<.����꾞�H?0'.>Y;�?���=9����Ķ>zؔ?�ZL�����ğ>s�?�t۾�n>`P�>�J����>	W���>s&E���':��@�=@?��iq^�bc>��Z>
d?��/��A��q^��D���y=�c&>��+>X��>��#�\W��7N�>��r>��*=��b����s�>z�?x�>���<�(?0�3?C��E���䜾5:ʾ�Iƾ�T>�ź�G���4��(����=�^4>L9�?�s�>�>���>)�E?����ᢎ>6�=?��>��>"�>͘?cɾ:�F?��Ѿu� ?�7�>"B���B=6�<�
4?��h>?&=�x�Qe�/�/?BA��0��>/��K?���$d�@=�=q��<��p��&����<�(G?Sc�?l��=�˾�h��]�?4A���蒾��=�A?���������V�R��>���>;=�>[+?�T>�o>�z�<kB��'6�>�5?�
�>�}z?�j�=�؆�b5�nF��f��<��Y��Y?Y�=���܀� !�/J?�:�>����*����%>!�@>��>�E��>�o�>\5ʾ9{޾���<:������w�> ϧ�dt>DΏ�sO=Ԙ�<��1?8��=��Z�=T�;2q�>-u��L�>�}��x=y��=oJQ�R��aG�s��{>��>�<���f$�T;�?�ޙ��QȾ��>��"�p�Q� �C�����,>�e>Z���}ξ18e�%���½��>>�������U?NM�҃=��*=�y���?T���@>ۿ�>?R�>
�j��ݹ���T��?�����{Ҿ;>�5?���5徘�g=1�3?ǲG>�j!��מ�Y�<�2=?A_�MOƾ	p�>	��>�諭�!'�*D����u��T=+ތ��lݽ@١�rޠ=㬆<�U���k ��$�>�Y>�����h�K�1?��\�:���}?��F>�V��?O�G��u��W��> ����о��?��>`���'F�*m/?�B�������>��>+u1���\��p�>F��۾`6V��l�?�g��5�辚0���`<	�?L�>�j���Y>���>f?�9����h����>�e��5ƾo��-!>D�>�������bf>=֔
><��e.�>�^*?!y'?p;Y>P�>�M�=$�?s�K>ݻ�><E?B�=U��?��_�a?٩�=�(�uٽ�� ?�3�,�>�>�Y�>Ж�>�ؘ=|����b?���>�������9�?����ƾ쳶<��G?:͝����>؋�?�E9u>�i��f��1�7?�?N>�����Ԯ8?�����G��;9��-����:>�@�?�&�>�<���9��ݓb����>�������=��?�^>V�>e����Q��|��>E�3?��V>fS|���:{?�=�oo?�6<�)i���� _�$���C����!��	�o>���5��<�)���[>�DE���==�mX>/�>�QJ�]1��:��i���:ݾ���Yg��1iq=��+�μ�`���\�>a]����>��>f� >�G9�ި`>�#D?�=(N�=��F<�����V������z��D��_�	>潓>���>)�>�(���W>�	�>�Z�^����x���^�\H1�Y��>66��v�=�x�=Ҋf> ��-�����>��t=�����<�.���,	>�⦾^���W�s>�˾@ͼ�t�>j�>{-U��^>Zv>0�?�¡�9���r����W>��_��`�<9~���	>��>Q�*� �>yδ>b{�;��<n�%>�-?���DF�+�=]�>�Gs>Zs�������>h:��.>�*�e������=�3h>�޳>/`ƽ�> ;���>SY�>wŽ����v}�9mN=����MG�>\i��L�ut�[]�>]�Y�Vn'���U��|>�&�=;7��~7����=y��;��#?s�Z>���>�2ŽFǽ��ؽH�L>!����2��y�$��J>p>��<�|��b�>�EB�d(8>\o	>�C��_=�J�ޤ������>���3��-?���Wټ���>MН>���[�����,����
/?���'e��m��f��>ިY�/4ս>ν���=�i`>7u���\�^=5A�J%P>n<>Y���t�n�?X��P�˽<3�="~>�#>K>%ͷ;԰����>��>�"�D�=?�c�W$Ͼ��?>�ۑ��9��LP>m�a>�0!�X���.;�>M�a>�d��s���٠�
>���c�=�>�.?)>M/�<�>睾ɶپfv6���(?��0=�@h��I5�w��+�>�)>�ߒ�����BX�>���t�>g
e>�+�5�����"]?���������l��'�zx�>�L�K �;PX�>\ �-/j���ҽ�g�=�+�� ƞ>�/�>5��B�>�U*>x)Ⱦ�S��H���2d�0�G�Ë2�<����=y��>�n=����µ>�	a>���<H�������tw�=�)?`Y�z�>�OU�����&������D A���>.TF�i�>xޖ=����)�=5e�=�b�'�1��y�Z�=�Dj����*8�=r] >�����s��	�N���=���=��Z�v�R=�{�>���>�wN����@:G>M6T>6)���+���1��p�Z>s��>J�=�|����V��>ؗ0=��r����n5>L{�=b�?�#"Q>���>c� �Dyg����a����˔�F��>iԭ=1m���wN�_p>�&?���~����F����><��=� ���z>B�/����V =�&>��<Ĝ��+]�	�3=t��>�02>v�߾�ǩ>vc!��p���A�>�4�Y�0> J)>q�W=�1���䕾��I����=Q��¾ӭ����>�����=���>9�X��ٽ��KѾ�������(>�㗾�g���B��S�r>LCO>.�̽@p=)��>��>�������>ўh>���>�}����>P�=�=��	��׽��0>=�d?�^����w>��
�P��M����=
f���aE����>hI�<�:>䩾���=��"�g0����P?� ��a&=y>��� ?�vo�<a�>T�>�/��䣼J�>p΄>RW>Yvѽ�%����=�ŗ���X��,�OFҾ0Ր����>E)�>��)>��۾�`>!E7=�X��Lr���=Poh>�$�>�����}�>���<d+���Ԋ>��ƾ��2��Z,<��>2���?����=�ܝ>b$�:�r�$Ȱ�7OJ>�	۾�v���W>R�f�	O�������Wv�3�>��>�a徊��=�?�3?�<־g^u��ۺ
fǽ�!�v��v!�=ĞE�J�̾��,�<�L>�Ͻ�����5�J>�� >q`�
(�t�p>3;Y>��1�T/�>3
P>�..>���=�'�������8b���=���	=-�H�E00?���N��������o>���>����T��|����H�>j��>s:����W�gx >:>�X=�a �6$��W��>���>�	�M���w>����"r���[��\�;�1�_%�Y/m��|t>�X<]�y���ý��W=�'>��l���>]��;�=��>���b�>�6��F�><s�V%H�(��=�Z��l>�&=nE�=�q:>�4
?v���r�Xs��ӷ>�#۾�]�x�;Ꮋ>�=�>�5L�0�9��<>
EJ��b�>0�4<��;l���䘽�b�<\V���<n�>���1�>��E�������!����/��u\������C\�>�N�>�0�>�Q�>�٩=4ӵ�z=� ��>@����"�����
�>�Q�>r4H��G���^>P�>s���$;
=AU>q�>Cmh�P�t�̘>ޖ>�]�Ւ��L���M	=����+��{v�=�؋���=~g�>{\��N�����>m��F�=���=!n;>������0�:��X��V����9�w+��8{)>e{�>NE�>&����q>��?���>ɂ>����o��l傾�N�#d� �>�Z�>jQ�>C)��W��>��!>Kk4>d�`�o/����K=ӏ+?�F���9>&%���;>/(.�p�����S�� a>Pe]=Q��>�*(>ju@��G>�UW>��l�a7|�4d0��\���=������>��>��9>D�>n�E>����b�����=-n��>���CĮ��;	>�H3>R9ὠ:�Z��>��>�g��S�>�!>+[">�/.��Y���埽u�>_p��nξ��ǻ�?H�U>�cv=}��>UP?I-=�>b��=�o��w��r�2�� j?Ò"��Ib�]6�>)	�=3o?r?�>�W��K�> �ټ7���&$(���4��0>�s>7��<1}��&e=�/�>���>U��!�<%�%�t�����;{���>�>}��>��p�>+�>5��>έ۽�g�'۽�%�>:R��Th= ���=�����A@��%�I��f����0�>�.>�
�> �<�n�>���>k.2�U����- �dL?�����Ō�}&�>��>�E=
O��树>Z��� 1'��Q��w�(<��>Z�>�	%����>�/I=*`�<Δ�<��>M�K�o�{Nn�-2u<>6#>W�����"qC:�p">�c>�a��#-?a�=�Ծ�u�>ت���y�L�x��)l>���𶮻�/>��>��n�U ���[�����>�J޾ݡ��/ý�I��lq>Ѐ�)�U���������j�;�
��>;=1o>mȽGE*=>����	>!�#>7
���Խ=Al>[b��8ԋ��@��7��=�0�<8gϾn���i�켱�>5W���=�?d?5>��Q��t��瞁>�Z>�8�<ێ��쯆>���=��!>g���� ؽ��>�]?<���9-���F���!�>3{�-$���»�8��>��n�BSJ����=���>�"��&
u�տ��V3>>���dƿ�>< g�>�q��b2�M!��Mo>��G��)����A>D�>�Qc�{e=��J����'>2sܾ�Fνs����޽�g�>7��>t���Rs=5��<\s�>�u���?���Ǿ"�>�A�=WLB>��Ѽ���>��>��S���E���-�8_�>!������ݽ҂�>���(J���)�>���m��=Ҿ�=]p=?��V<J>R�<{��=ݶ޽�u��t)?A���4�	>�U�>T���Í�>W%9�Q�����*>�X�>���=��ؽݣ��
q�>�ӽ����t��B��>T��>	�t>�,��@�sӹ��ќ�L3��ČQ>�����ʾ����d�>r�e�lg����ý�o�>Y�>Ў�ʴ@�gɱ�*;��ˢ�������Ͼ͆��TgԾ�f7��_�>4u�=m�:��I�)>���=B=�&ľ�R�Y�<<�E$?�u	=~�/>�a�=`:?�i><޽eߟ=� >�G�>�6@�	�.9����?�E>2�����ھҐ�>���=QI�`6+�s;s�R�����f���t�]��
m�'Ó��Ꞿ��@��a>M򋽔S�=�I�wT�>bn>�ܒ��Ϝ>b>�>��?yj�?ӑ
?�>��9?���>5�>��?"?�)?��?�|��.���YC�$�o=t]�=���>|��=�9?�Y+>mG/>��>�	<�6�h�e<$��=��	��Շ>1��:+;���>ꫩ��h=?�쾹�y��{>h��=(��6��>^Ɍ=E�>��>)t�>��=�U�Μ�>N�~?�kʾ�}A�->�=��o>ƈ�(���"�ϗ?�j��q�/=�|)�AT�>ç>3�>��>�{*>sX�=�߽���=��
>�YA=�)>Q�?��>Rs+?��>��>J,
?��N]�;�;�?z����=�E�>�M?r����=�>��#?�3��"^��WP0����<���>�#?k��=	�>��E���7��r�<t����'����ڨ�= ��E�,��ϸ��V�>y� =�)�>�G
?R���l��K���� ?3N��1������G��=gfJ=��zj�=�k>=��=����+U�������5���;�3�ѾҠ��;������>/1߾)79��`˾H�cZ�����������<.�T ������;��fi��M6��
��Vww�
�)�>��K����
�!a��ѿ�>v�߽��:����A�ř�+�=�C���rؾ�N?��>?�6ټKlu��#�C�>�<�Vnﾵ>	���>�O��<�<~C���q�J�I��� �H�@BI�t%��;��=D��=�D�<�>���>������>º?�ڳ>��
>S��>���>��H�;*־��?��M����=�<'��p<>(A�*o�>/T>�j��۟�h�>G׳=�<��:?Næ>�Y��k����>3ٛ>�kƽ�	�^�%?z+0>�+?�@>��O>%?X�ľ����.?hԋ>�Ge��D��'B߾��q���J��n>���s�X����'�=��=�f�>�J�N(���﻾(�?�9L��-!>��>9�
?�~�v�>п?cr&>�& ���[��6 ?�%>L7��^���)�|c�=Y���$�*�*J={��(,m�AWk������X�ëm����^k��b>���?��>�X_�m�>�{>�ş���L�-��G]J='yA?��^��>��<b@:>Ѹ��������ڡ�>�P�?Cc�������_���>�����_Q=%�Z>c#�>�%���Ǆ�v/���K�>Pǅ>c8�=�H�	���v=����?�;��􇞾�սmu>`DG?W�R�>�%��e�v��>S��$#>���=�#>�Щ������e�}��>����ZW�7)s�D�I���L���L�w��6L���QԾ���>��>#�ƽ�?�?�9T�����Xp�KY�>����]ؾt�!?�N�>`�i>�O�>��?r����r	�q�9�F{����=	Z:?*p�VD׽�S���ြ0Cͻ����&'	=���=;!?O����m=�?->��?��]
�;��?�d�=v|�=��>	Թ>��=sa�<+,=�Z�=4��.r[<b𩾘te��!?p�>$�S?���>$N�?�E3��"�>�?p�M=a�����ʽ���>@�->Ҙ�>v�(>#�&����?^�(>ޞ��5�><���#>�ǖ>Q�ʾ�n�=q��>��f�oL=�s�?� ���k{<�r?^�?��	���g<�fN?�����ѻ>w򋽜~�>��=��>?_f>0��>N���0��:��.�W�;�9>Ñ,��Q��*�|T�>o��3�N;�����(�=kN�=������<<�>�������<(����w��Հ���?F�G?-@��飲=�Ȍ>�3?{R���>�F��3?5�>�
��6#*>�q=�͝�HS>j�=s��>�������[	�0"=O��&����0��Lټ<%���~D�0��'���5�x=[=#a��qC����>��F��a��}���IN=OZ�dj9���q������	v�����fν���jX�>\�?�d����!�ݽ�]n=@����J��v��P�d�]?�r�>�������=�x�9�o��A =�<!1f>�Ҿ�j��j/��[��&�> *��ݾ�ž���G�E?���>z�ξ\�E��Q1ϼ��,>��C�X��>3�l=�g�=Ml7=���>Me��T���5�ü��>�?��>@o�����>,,<#{�J������>�6�������;$r�>��=^o̾a�=i8\���Je�p�>�{�|g��@o�>3{A�]�-�.���9叾�jO������s��A����ξ�.�>F��U
�WD�>U�
>��M��w4���=�\>��=�����B?���>���>qf��ג`?�p�� 1����V
�>��ľyn8�!�_����=��>�������>����?c�$Ś>�(�>�%¾���C3?m\��ǽ-�����ż>*g>�=<-�W���=9=þL��H�r�L��[>�D��*��W���=��>�Y?u���K�8��dL?\��=ۓ���<����:��>�=J?3��>�t=z\?�0�?.�8��GJ>���=��E>yT[�~��=�:4>|��=  侠g�>�� ?��=)��=��W�->:kW?�0���_�
k^����=Bz̾9�?���!��?V�
���k=�X���r?rX=�[">2sx�/�K>n�<�;����>���>V3�<�f;�aM�vrC?τ">��e=h�����>"=��}=\��=�{>O�=ǈ-���ּhOQ�E?�O�2E�=)��>�u�>��/?u'w�����x	�>;
�>�\>ӳ�>�ؙ>�X>d��>�U���l7>����k�>J)>D�V?�4�<#��>h�>Pس��Q&:��z=D���c=��ʥ)?�7����7>�1�>���q����0�Ӟ2����b!�>�w����o��=8��?Z*�����Q���5h>�C���zI�������=��¾
;���]�>�ǿ�u]K?��Ӄ?[\��`�>v�??��H��>�S:><w�=�<W͊��p���4�>W�?2}�>��
��[�=-	�?0up?gP|��Z��|�>���=�t�>��v����>:x�=3Ϳ>*.i>��=2�½;�k�$h8;eD�>�ʽ�Г��=�H�>�2�q%;�b�Gf�>���1���ç>i��1|����="���@����~��.�>�����Ę�h*�=�zc�/[��/�>j��򊓾1x���j��7ݾQ|�PÌ�磓�To,�K��=�O<��>51����ӽ��۽+h�¸R��Ǧ��nǾ(�@�WX��ύ?9?���C��>��>�/�=��˾�>GP5��=?)⽦/Ƚ����k� ��;��}pS��[��g�?8|��p�<F���+�H?c'�Q��<���>�=+n"�򤚾�?FSY>VҒ=�_���,��h���qd#=ԭG��94�WB���F�?B}�����8��m��^P���+�Ұ=L�4<���釾�����@��[�½k%�n��>�
���<�u�§�<C����������0>�G���m�����v�?�H��o��Ƚ��pg�>|!��٣��p����b������~��ۡ>o��>��1>u>��r��2c>�����2���,���>(79=s�;�x>�Fr>�QW�Q�_��~�>͹?��>dݚ='�=j\�>��4>�=^$	?�'�>��>Q�;?}�c>'�M?�?n�'>B/>��\��%׾��K�����^�>�� ?ɇ>���>�#)=�GD=�JX�0y?B{��������<} վ�޾���<�Ϳ��=��]�^D��H�4'���Խ	[��5,����N��c����þ9`t���z�����U��އ>�ч>ݡ�>s{5��oc>ZE���e�;ְ��������0�����?�d�� ��̛��,�>`-?��ƾ�V��Gd�2A��|n־��w�@��֖��`{����/��⟾a{�²�>_��y6>_��� >ܡ�K�\�Ĭ�=��K����x�ۮ�8�[��n߾hX������}�>c���c>�֬>�i�>%w}>V(v?1|x�_u	?ZT�=�:?���?AN4?��	�$�>t `>��>�|�>�6�\��>��?���>�ѵ���>�$$?�Xr?��)>pN�>��O�4����d˾��=Y� ?�p��ȁ?q��>RN?8d�"�g<2?��>0޾�ҽ70#���>�ő�:W0>�g)� �>���>�t>�9�=��!=�h�>\��>N_�=¢����X>�f?\a��g��y���?�=^��]V?z\v�-no?m��>]�+?X�I�ºS>'�s?Yp>p��0~>>���ʃ>�&>���>�_�>ت��^y~>Q�����q9}=N�>�����J�<7�I?eO��5�=��=��-ս�j��R���\{>|�ƾ(��y �C[�=7���t��!���(��=#2
�&��>I�w��Q����=�`?�h����C=��C>��>f��;/<��QY��"D?��\�|���'�1?�{��ke=��>&���Yo>��#�q�ɾ7�{�5�>�`C�Y�^��ԓ��8�>ʭ��2�>��&�1_x>����yǾcUV��`ͽ������[�~=J���0���D�G��E��^X}�늌�I#��N%?cݾ!L�J�$>[�
��l����T��i��q�<��=G�8>\eN��>�c�=��>�3����J�:*g�*�3��]��?�A?�<���>}`=B�?�~ �N캽9�	?�)>�Ɓ��p��ϧ=�o�=��ξ1W�>_0�LM<?f�>�ު>�>�u�=8tf=z�i���=�l�j���c0���,�4���t>/*>��9���M>�d�=�ʋ>���=^��<����uF��6?�P>J�ܾl۽���O�/]t>��?\>�-wZ>���>V�q�����5Ϻ�WH�>�>���$X�=5��l##��J?��U��V �6���Q�'�>��2�w��>�F;��{?�~�>�	>����1G?���>�%�>��ȡݼ;H>`�$�����>����Wm[� ���¶�>4>_��ڴ����>Z]<>Q�=��R�a�۾�0-��=ľζ����>C��(_��#�'����=�&�>ߋ��7+��V�>�+~=��<�6?�I�>�6���6a>wÖ>��?�z&>��>p� >)�➳����>�I�>���ފٽ!����>�������>ߡ��=���=�F#�&��Z��2�N=DAɾ:�	��X=�I�>o4�=i�(=f%T>z��>u��5oӽ���;�����c����mU��t�=�>�	�x���c�>23_>������Mm���4���+=���=W�z����>�v�=��<��^���=�
�>��=�n�Ω���?
�ދV=y��>T�?EKc>�������r�ｼ�O��ͻ<�Ց��?L��M�i?����2��9?��?�>+S>�]�>�˙�8>8H�<O�A?4�>��5?���=�k>��?��>��>!��=����R�#>]Rq?���<+����R��_�w�&Y>>�]�=�ch>1]?��۾]��>���>���>��>"�?�_�س�>�RO>�3(?C\�>�^>���=�n�>�	�;�}H?�M�����Θ�>.��'E���hʾ�꼾?b龊q#��~K����=��X�10?s�����8?���=UoL>���>�� ?`o=�腽3��>��?�!2?.�?7�>��k>�qP>�X��٦�>�K���<�8�>��I=���2�R���>@F�=�3��,����%�xA���־K��������=�9�>�Q>��<����>O8?���H�>u絽��������JD�!^/�h��=��M�+ˁ�;�$�,Ï>M���=�&�ׇ�<�=C�I��y1>�1$��{=��ާ��?T�a>�3E=�>n'ս#`���¹����>ā��H��#�����Ⱦ �<��1>��>[f?����Y��='b$����y��=�!4>�0�����޾������;�=ɞ�;�*g���0���Vf�w:�7&�>��W��c�Y0��R�=H�ž��8�z�>�.�>&Ʌ�	��>�G�u��+������b=�˨�S!?�/U>�"�TM�k�[���5>��Q��T
�d�=,�#��sA=%iu�.�>^?�Ę�,�>Q�l��?d����L޾r0��J?����(���M�c
?yy�>879>9Gi>s��[���1���t�Jo��	��>dE�0�� ��;B>&���
���K�O�l�x�}�~��:�"?_�c�<)�>���>]d>tn�����>P����!N>�+�{�*=]�o>�U�<-����>��>�4R?�u�=�R\> kD<0�x?��-��=��	?�9>�/羍
�0����9?f��[Ű<�V;��X?�Z?�S��C�K>��?�J�><����>lV�E�?\ʾ�����'���Mg<��˾��.���>ޓ,>�?�;*��=�К>�g�>:�0�<�>�u>���7�=�5��ľa�b�q���Q����>�蹼��>�����Z?av�>��H>�"w��?���>�z->��޾z�M?_s?��?f�}�L�>'�`��� �> ��9������?�~D�<�~�(���"�v` >�<��x��I�s���X?�D4�/��>Ԉ�>ꣂ>8--�>��>꯭>��"������.�<GT>�̇�g�>0�>��?aӾ7s�=�q��g�9?i���HP>��>^��>5}ƾ���>8[ξ��>�V�=��<q_!>�
�>�F����?��}?b���K�3>���=�z>O�,��T����'3i>��=�?�O:?�0?��>��m�xJ���4Z�ϟ�>�*6>�`ƾ�?�̣�>B�>6 ���;I�CY"�'���b�,�5�����">��u>DZ�>
5�>�5�W��>'�>8>���S�> x�?�w=nQ���R@�&l�>e���Ò>��>!E�<=PP�>2�?�@�.m�>.-S>�J�?(a�>� ��AO����"�Z�W�۾�:�?��=�A��	�>	n��)?���=��8>̜=@&#?ƚ=�󽵴r>1�}?��?�a?2]��غ�>>L�a�/��Im�c�>G��=(��;����>�y�=�V����=���>M���}Y��'p?��>t�=6Q��y ?�����=���P'�A�d= �Ǿ���=*�n��`��������9F��)׽�Ɏ�l�A�������>��!��r�&���+k>-r���A?��%�Ţ��^+��=�KT�m��=�о�P��!��GI�>����^�׼��܏�>�Ԛ�S����>�?~>�|����<��}@�=�٦=R�=��e2�B�
>��a>���A�?%Թ=�O1?7�ھ����s����;U;?b�D�й6>-d���>�<�2��V��S/g�v�۾��
�������=Cꋾȟ���'�e�6�s��>Ǜ*��dG>�uG��'?���o�̽C�,�����o�ho���^=�殾5<��##�Si��&��=w�|�xK���ka>mj���؂�Y�<?ךx�H�ؾe�o<���uB>c��2#������-r2?�ھ�nY��26��?]U��d�=m�o=�2���씿�;�����.��������$�����tϻ>��>X?���>�0�=F>Ro�=>*`�>� g>�ǡ>�m�=`H3�A�>��
?�
�>��ڼ�s���Z�>�>]���Q�7;]�5����?�Ɗ>(� �h��=�>�������*�K��>t㏽��=<ZH���>�f��Yƾ�����=Ό���2�)���0�=���9�����v*�od=�V�����{ ������=Pf^��_>��<�:U�;��>�b�>�Q��U���"�m�>��=`�H?i]>8_ �N@���!���>��>��۾�#?���~���%m�6.����%�M��>َ�=��
>�C%>�*?�^��q����$,��>��A�,ȅ�ev~��-h��Q�nG=*_���K?r�>�B��>n?8y7?F"���>�6n>��C?YP�/~>���>2P$?I�ӽ��3?���>>�> �>��)?|��>�R=��x>�}o>'��>}	�j��=�6z�.���<�*]%>��ž�������>�������H�4?�j?*оK�#����>���>00�KuZ�h���Q���{|�7o�=W����;��`>���>��)?�ξu���ž��@?�(��qޫ��V��|'>���C��=�� ?#l����?G�&>�[>��E?ȥ�>vǅ�Eڠ>��}?�$>�=� �3�>�H�C47�Y=@>�p>`�U��|u>Ga�>G � ��iۙ>��=
���:�����>���(���p��;P=+���&~����R���N�+8M���&�;c�=�0:�66��������>c��>�<�!Â>R�>�Q?XT���o�C������.�35�>����������5S�.�=��˼�
��b�>�Q���%>iGͻ��=󄙾���>rD�=�
��tU>/٠��U�S���D�>Yܽ�C�����=:�����=[�_�+r�!Tʾ�����=0�F�����a����E�>����/��O�a�T>���]�<Y�ǽ��>.�>�T=5aa>��BՀ=���v��>t��ư��'�r��= ���p�d�jU��o�龛�>��_�j��=z��>L)?=�+�������=C��>a���T���r�=tq�&�>B�/>p�6>��R?�����>_�D?���>�P���T�=Nb?f|M��k����}�ž �*�Đ]>,ξt6���?>�`.�a-�=�Is>Q@�>D]��J����u=�>��=�����\����=jVo>;2�>��>{@�ذ�>��>��s��Dn>�>rx���>fn0��
��྾��>M��<5>��*,����YM?Y=�:N>�E�@H?j�>��>��>�(�罉�>�
h?,��Yݬ>P�b=��O>D`���G�>�'$>��=�8;��*r��Ջ�E�N>�aվ�]�>ҾB�H>R"Խ�l>�?V>�IS��[7=��<<�)��.�=̏7?B�?X ��G^��/�>��t>�\��q�2�;>Ri��|sV�r�=}}K< �=&ϼ\�z<���Br�c�(?q�}=얨=t���*d�>���=�����(�>@�?=��ﾜؾ׍���i+5��>�1�>#��>oK���?]�F?%z�;�;�6�ýeh����J>�= �k>V�<B�(�ݾu�Y>@Y>���tqؾ������l���K>M�#�J쾞gd��>�1n�8>�j>�6�>�.��]���L�=�x�;Sc4>}�$>��>u�>臤=X+?���>�������h���Wо놁�z�d��N/�=�=|i?��>Z�,?f �>$L-?{������>h����.=�)K?�b�>�p>�矾TC?��s>��>5ٽ:��>"�>S�o?<!G�یd>�>���|_��m>{�Ѿ0���qj;@^�>q �0����>'��>(p?��0?^Z?_��ߢ+?�a�>G�>��>�#v>T�!?ǉ�@U�>|N�>nvw>�a��zt��{!�F�k����=��j�	��=�\4��EY>j�>U,��-�L�?Ȳ�>b�>[���.�>I�2>�1?�J�4Zh>�0=��U<ڃ;>�PF���*�*�v>��?iK	�gΉ��ʾaZ�>�C!��lC���þ��>F��=X��=��G>P�ʽ��?x�>�ԽXƽ���>=ҝ>s�6��[�<L�=i����N�c>i��>����
xe�������<��s�u��K�����>E���5^>�Y���PC?��>�|Z=�7L>��p=��L��Q���]>��� s�>��?D��<:�p�"��.�w>�<��8�#��=���M�= ���\P¾ˏ;�љ> [o�	M�?`Ծ��hks�h�i�.�7��u�+��>�CL?`J?_֙�fz>�8�>!��>Ľ���ց���F=��5���#�I���h�>'츾E�k��	!�mB?�B&>1x���,>N�=Ɗ�Z<��������<6�Z���2iF>�c�<q��>Ll?��������{>m�ﾽ��66�U��`~ƾ���>�x�4[<|����S[?5ʾ6m��@3��L>���>������k���>t���M =b�/�m�H�'��>�TX>���{Ka����O��=����N-���+ݾK¾6!Ծ'����|�=�r8>j��S_1?R����=r�?w?�)�)��<�I?M�!>�Z��K���X>�J�={���J�=��>��M>�-���=tG�>��?��^:�~P̽���>���y���8��gٽ}��=K# ��IM��V�>U�V?�̷>C遾��>���>�U>C��<�D�2 ����NӾ&|>�����Uys�X��>f��>�"�5�=��>�F>w*�ͺ�=�r��B^��.�꾑��=�w�.P��x\Ž���}�8?XS�=�L>d��2�B?��>��.?��X�kj�=��7>¦�?Y\W��=�|;>o
2>�����=��> ��	�.þaf���~��@�{8�=t�A�)����uW��u�>nh��Yp\�6!'?�Jh=L��=�׆>2�>��վX���?�A�>���A��^>0�={q����>�҅>���>��\>�S�$�0��Ζ>�# �	#��H9�=���>\ɕ�0F�=�f>��?�VA�~�Z>�|�=��>�����(��()>��Z?^�_=fwu>�-?�ܾ��)��|?8 �>O�󋁾�9[��L�=j҂=_h�=� �>���E�8{e>�Jb>%p#��s���.�<��:�Ӌؽ��_=���g㧾�Q�=�? ?���>u�(?��^�zH>���=�&3?a� �ǈ��w���,}�>6׭��{��2�>u
K��%��j?pB?�����D�!��>�>_�=�޽�ӆ>B�n���]�Hf;���>�����=B7��R��(�Z���I�7�?��~>E��>�1Ӿp ?�N>7 ?������>ދp<�S>�ѧ� |�=D�������
�!?�?Dh�����k ?��=�>�ȼa��=����H�c>���`����g>��@?�ʾǩz��"˾<$�>�����b��H%��N�>K̾љ��ߑ����&��a>1>�����*�<�3;c>�C޾��e�~���B?IЌ>�r=��*>@��>Eݞ�ȏ��
���ݼ�(�6nS��Q����,?���>���&N�<�?��?�E�=*� >���=����y��<0:T?p�v�D�>�����>9L�=�u�>H5���7����=�U=?�����=��ｫ�H=�O>>єA�*����|Y>�J?D$�⦿����R��>�*���qQ�Z�
���>츤�)�.���޽sv}>u����'E?>�?�ƾ�N	��P���"�>���[٨�J�~�n&>3�����
��4-�oU�=��>)l�D�����˚ܾvB5�2?i�s=����u� �<?�+��~lp�Ё9?.#���b>��+��G����6��й>
-�Iu�W���o��>��Ƚ��Ž��R��?�M�<}��>;�~>�3M?��=D�>�<?��Q?�v>��!>w`�>����B���+X>�Y˾]�x���k��ֱ����>�w?__6>�6?V?��?$Ӎ��iQ�X�L����潝�;c��.D��nQ=o���犾�������B<�x�R=���3�>Y��Lپ��cǃ>�\����&yu�9�;������%B�Fũ��h�����H�d����Z�h��a&�R�|J>�ZB?ǜ9>}�t�ו6>4�<�s?�g��f?D�1?�V">���>��>�r���콗(?��-�
41�H�T?�㾔b�������g�b2d?�i�<� ?������<2�G��e�Z���,�T?�u��|J#��š��!W�-��GHӽ�u���@�Qv>�DS<LFi>�B?
��?|�>?[�?*�A?q�&?Q��=����?�8?���>�y?C3�=M�-?Qu�>&qj��r?�?���>�
>��=�">WࢾP�	�� #���B�Ʉ輗�����>
�7��Y>鹼>���O0A��-�}>��9?@�m�b����3>�ȾJ!�<<m; ��~���>�@���=C�����=�!=OO�>s�*�V3�<��꾀.
�t����
>>Zz>�/�>(�?y�@?��>v�?�¬���>1�ľߪ�>�:?@�o< G����?j��=�~�;���l��=�pӽ��=�ظ>l�X�6??��I?�o�=�E(��Q>�j��_�:��f�r�ѽGq��4ㇾ���&(3�ݣ߾�`f;i�3�t=���\���x�?d�"�_4��?�=q��>c��=Gg=þ==>>����ת�.C�=�lZ>�Ӻ��0��I���?k���o:����D>��>��#�ig���!��,�W�D�.�2��If�VK�?�＾'c.?����|ɿ�'���˾:�!� M���ᾠ�%<�"����:>D�C��M��ƈ�����,w0�!�l�m�C��nE?2	��	J	���ʺ�y�<_B�2o�XN#�+�z
d?�#E��>�	^:?�;���V3?��>�~W���?>k���z���w\�1�ƽ᮳>Zq�>x�>�k���9û���>�ݲ��������г>�A?#�B��ve�La'>|�C>�M�>�i�=_�z>��>Ń?bV>�?�¾֟򽚇'�d���_,>$��3�>W�=�Q�h��HxB�����3��=yj�K�6�>&�?����b��q׾������>׬��ŵ>:�8?u�>�x��PL>CC+>��O>�oO�
��>��]����Kr>M�)�Ҿڽ���>P�����P�Ӱ߾V�#�"�پ�U���nr���D*?D�:>�S<���'?(�(?��>�(��4:?���m�k����>�?u>��>�
������"��e���վn���"�<(��=*	����<᳈���Ⱦ�Z"={��=�^>�H�?�f>h6%?I:p?qf�d *?�9<�(�>��^����;�Z>|>���(���_�	�� ��X���Z�s��˪��W?�)S�?R��ξ�O�{]>���=�p
>jW2?X��>�)Y?�=o �`�f�����o>>oYj����>�q
>D�>*]4��7ؼ��x=��켂���B2���n��𫿾�w������n5�>66�x%�cJ-?�T<>{�`?�+>ƚ$�#�=v�JŚ��6��*�=q��=����mS����7W�b�(?����K-�� �ķ켾��>��U���>�S?�O?�/k>kT�>.^�>S!n���'��2�f���܄>�&=8Cp>0]	?Hmz>H;?Z���H>���?>�=[�=)�<�&u�J��>�<�>�>e���9L?O�`?LAF=n8��RA�>�Q"��(<1�=?��c>W,�x����*����J�;��$?��?�|�>�I�?Kꗾ���=��>�J�nn?���>����N8?�����?/��>*���M��>����C�:��/
=�d�uf>�=6��,2�n�3��*(�+Q=�X#? �1��܌>Ql�=�.}>Y���z> 1H?�����?��>�0=�ܽ�(>>�?x���`�>��
�Q+c�&�=��������f�6ؚ>���>��i��ս�I�=�?f>n��.!>�>9 �>!P	�0�9>*d��V�7?��6>��U?���=��Y�\ʾ<y4�$f2����Jv�<���9�˾A(O�D�Խ��׾�h"�����?u��M�羚9���ɮ>�A� �>	e�>��F��6��bp���D�>S̾��?�=����	��HJ���E>���f����7>kj�>�A���>�]���>'���q���V���%��ê<�g����?�$
����>�2��נ����ľ4�>v��=���j�>;}��X'B���'�����-?�3��c�?@������I�ҽ�?��]">�M�>\>�=��漈�u?C�9?uY>It*?�-���������Y���������>i���ڧ>�����ݾ��= ����Eg?��ᾚBf�S�|<>dv?��c���þ����B�??����a>=>�dt>^d���¾�7ž�<�S��t�<��$�5�N��VнY�;>Vd��y�ɾ������"	���e�q�L�:������h>c��>?�
�`%.?^o��=r��]@�d��>�Ə��2A�C �>�j? ��=����~��޽4?�M?�ૼw/�=�EW>x%$����<QB9��\!>O�^?񑬾)���ͻg%���qF��\�s>7¾��`?���=��V�ۆ>U��>��>�n�"�3�/���"��K��Q�%��T��_��� o'�J��>�r����>�a��g�?�c>���>�H=�Q���l�� �	��� ���I8��]��y�	>���>�*��E�>�^:��w?�F?��=hQ��g�;?���>R��=e�+�s ?��=	�-=͹⽑����;���Q�������;�]�nx�����YhϾU�������}о�_��&=t��9�=Mי�K{���]?�T��b���`=Q��m�=� �>P����}�=�E?N��>��>��L<:n?W�">yה�WVþ�?����7d�eM=�ϼ-�??��ʾ��>>���>��?�,�>��?^�B>z-)?�^W?w�>kJ�?�.�='�𶞽W�h<��h=�&
?�N@<���=H�o>��>Í>���J�>��Q�F��=��%��d�?��J��?�S�	�*�c��pY��$T��?U����ܟ��lվ�R*>_Xоf�T>��7���>�}�>)��>'��ҹ=�ƾ<��=���	�><�>G>��=a�I>���=*�����>&t?rE�>�$���>�ºuE��m��/�ž𼫾az>�WS��1\�H�>4��;^Y->�;���pH>$�I?$�?����P?�̓>�U>\Zf�蛃>���|~̾�0`�.C?��>[X�%���jƣ�*��>���n>�Re�>GQb>��u������1��E.��s@@>� �l3>�����Ԍ>��,�����1+>��5?�7������e�����Ǿ4E���d>K� ���:�9�ӾEpo����>���F��>k?7��Wi����3>O�"��&>�ZK>�\"���>p.�n��>g�>���������=G�>a4�KE�<_X6>���>	޾5�������Z�E�}��=E�i=�&?�I��k��Y�?�}'?!�'?V{`��C��	&>�A��x����>�dB>�R=��>�Mw�|�ֽ�Y���Z>��Q�Ii���H>x��> ��-��P���B�>�*p�.�;���>Ϡ�>̷C�]��>53'�'*>UW����:��(=��?ז������mG���Ͼ����k= K�>�o6����t�>��տ�=�$��O��d��>���R�!�C?ػ��)�>��@>t�G�9�>�����P�>>"�J>:���Ñ�����<֥>�9g��>>�a�<��>T 5�{��w��>?��>U��>�"�>�|�>L��>^qR��d�Y�=IY�9�%=��L>᜽f^��{>��I���`�>=`F��b>�c|��6�?���;����u�>Fri><� �^9q����H>+��2}��D��]A�>1WV�����|��",]>���<w6T�%���=�?�:x���ʾ剺�k9�ԊI���ݽ�6�����7cb����۬ؾ1��>ˠ&�֬�>룡>�%o>`G���J=aq4��`+?p��<��*>�{[?y_2?xN ?B���.��>/���*?f�T��c>Ҫɾ��]z�d}�>��˾��>B<sV5�j%�>x܌���=�K׾������R���E/��X5>�D��5a�M�B>EH�>�3��:��N�6��ڄ�3.P=CX�>��>?rm�>|H�=���G�?'/�>�>y�g>�H#?���<� �,�?��>�M?flc?۸�>�6?�A{">8�=�:˾�_c=�ȍ>�@��-7?��Y�8�J��L�=J�u��o�>�L�z>`�@����>(�J�doE>�_J�z;o�#��x��Yw?-#�>F�t�'�"�=}�=�aݾ�¾yh�>Sj?��Խ��ң(��Os>8ם�;��>֐p�AHD?�ƞ�@]������
?,˶>!m�>��??�\L>n�/>��=��=�g>���̋��9�,���(?�lu>;�E=��T��?F�/>�?z7�>�3�<����L���>`$���Θ����>�g?
H=g��\]��%��=X�.��3�������6����>D�ƾ�X�=<d���>wٞ�Zy)��Li�/�9=}�>�V��K�%>��?�	ؽ�Z�iN��`������>�Z�z�?g�"��E��0��c�>��(>�\�>���>�>�>��I?"x���f�>z�T��Ã��
W������߾w��.ߦ>D��=�_��+�=v>e;��(ڒ>)�U������A�Rn_>t�	���ľci����=��u�al��l�>^��>V6��F�m�ᾂY��c]8?���*\�>��-5�>�m꽜Q�č�_7?)6�?�������7@C�#"��,��IlE>
���G����2>���>0]�P:d���:>hrw>po��S'�(v?�+�>k�������a8>��?�N?k>��?�ʷ>���=�����>o"��J�M�g}��&��?�`�O�f2�>�ս ��>�띾'��LH��(�>C�N���Ѿm?�g?�?��$h���>S�?��>�Y>{I?ץ�>M�q�W�J>�A̾|�n�/'�j[V?����[�>��>]�U��d���|q��\�s��8ƽ����6�>gh>o�?ҭ{��A?⣽�=���=X&�?�ܭ>����덾0� ?�	=�"P�>�q�ő�̻񾊁���Ղ����-��$>+�Ǿs�> m�?���>�E>#B�>Ja�s?��>C�f?�ݷ>�� �����@��?�Q�;��H����X��>q��>O���i�N�����#
c���?�nb�	NZ>X��>��ʽ9����>35?��s���Ͼ��u>�B���=?]F�>��y>����yk=�e9>�Y���y�UE$?���>W2��rϾ���>bR�>b�=?���[�=���>_�̿�����I?B�=�v->T< ����>��u�ھ��.<�?5�?�s�H�߾R`�>쳽�E��v��=�;��j�N�(��:�>JcF��l
��>?" ?�gQ�ML6���P�g?�i�>o��>q�?����#�;$�;��F��_6 ?m�=-v�>ioɾܥ�>� =�ҷ>� .�H��>��?�᧾�%2=�-��vk?<6X?Q�&?g����?F^Խl@�>��Z���P?���>��<i�����?g�V�ܶK>�	�3#v��?��|�=5S.>��N>��l=mx����>Z�Y?,�j?��\��� ?{�>�ۖ�J�9?�K��6U>�%�>���>��,�e6�>?�S�7��>[���>L�>��E��ȼ�C�,�O�f+0?�g��jg?>�?*�8>c|��Y�=N
�>�2?C����M?�?Q>�q�^ˈ��F�=��>LΗ>��=��12���>><~�>Q��4���KR�}o�>	���t�����>�f?��u<:H����>Ʒ��B?�,�=䓾to�a�B=���=��L�Ņ*>=έ>.;9??Q��I���g���߼��u��0�U�󾃲&�[������S6��T>�_�"U>�@,?`�B?dw�	�J�,��>%1�='����e>VD�R�@=_Q?�%���r���!)�& �?ɳ�Ͽy�/Q$�S0E>���>��=�&��^���sȾ?����MW�ro��ڔo������=>~(m�mq�=Q��>)C�>|E��`1>��C=��>FV����5�;�o�?F��4矾�W��p�,<Y��7u�;#]H>�1(?��6��Ӿ���>G@�=�����?l��>K[�>>�˾�>^��3��=s�þ�sr�}�)�ɲ�����%[��GԽ�D�=[���6��?@��T��`=�����>�B0�:��>bB�>��?ي�4�{r��~��m/���K"?tG�V���gB��}Ҿک�o�X�z���l�>�]�g����F�>��|?]�콫F��><[x���4>�� ?�	�>��G?�s
?�ڽ�P ��**��?�B��M4���I�9��>�u�>S�����o��?Y��>��h�J��<]*O��>s�o,�j�=��ͽ�8P>Ȋ��zލ���
?���>��*�g�h�k����Z�=�>��!?3��>3����A7>��=�K{>o�>����>�p{<?$�>'�:�����=7�<�=��s?�m�>������H�a��s>��.d�>�*>�?�X�N����	3�a�F���z�>)�^�8?׳�>�7?�P�Wn�>�`�[*�>%@+����?[� ># ���fW0?6ل��?�:#�ɈJ�W
`��>ӾOm�
8����=zu�>���3m�=���>���]���Ͼ@��sI�>��><�ڊ���`�p �>�^�=b&]�U���&i$?�Y^>��8��&_��Zi>��> =P<��F�?i�3>���F�!��$�>�҄�8&��D&?�>�'�/2��+����� ?X��>��i>:��?5��>��?���>M�?	��>߶�>�	׼�wu�">�Y&��-a���I�*��9~���>��>��Z�>�M&?��=�1�ܢ�f[v���8>��q���3>��>">f>[����� �PQ7�軉�/־d�ƾ�8E��ޅ>�D'?6�v �>�j�U�>:bB��=?���=�ձ>#�Ë�$vG��'�>�m�<��$?�]y>�>����تe>&j�=n�2�ap���=\?�K�>0� ?e�u��멯�u릾����a}�>���>�|O>s'����>)�?��>G�
�6OH?��%>��g��@��U�.>��>�=��ν]�3>IR5���򽔸�?��w>t{��׾�%2?�a?�y���E���-0>2l<�V`R�Y�>��:�	x��r%���ְ>�A�R)��%��/�=y^B�b�̾0�l>�
�>~S��\��↩<M�(�)�վ�~��~�=�Y���-�8f�>��_����(�?e�?���$F���>���=`�t��N������Н=1Y��}���+�!?}?$��~D��6?�c�>��+�B>T�DL�>�f>A�ؾM�L<�>��>f�>jQ�/�?X��>� Q> �<���?� �B��f���"�S#%�]�=|y�=���[��ì��b�{>�觽~�$�(lT��v�>�_��yL�T��>i�>�1���"�f� �Y��>v1���,��`�����>R���G� �u���#� >qP/�1�ž�4�� �>�0�g�7�6u(�a@Z�_�_�h����>N�I��i=xu��e�>Gb'=c�>�֍�� �Sq�>C���W�����?|�>�$!�x��m���>%�Y�#M����;h��>/Zݿ;?F��F<�-�>v�F>rn�l�N>�/?��_?3�?dzd?�	��MϽ$Ox>���؊�>����O^���n>3N>��A�ت�>U�ɽs
?��U?���>9*� 0��<�*�Xg:�ꣾ��>�;=�I��=�=zCE���Ⱦ	)>�Cݾ��?k�?���
����g=�=8q,�~]���J���<Η��Ҿ��=���r���K�="Z�����冡�G)���Q���l>��>����{BA�V�?�V��H�k>S�>��)?�V�N,;�����q����#?�6b?�$�>Z���P�
?�pоФ�z;�(?��1����>|����/�>Q	��CD��1�>���>NG�|��>0�M��L�>U�!����u�>L����䶾G��=*�=�L/=�\;����kE�85��y��>0q[���}=�5>9�>�|A?>��{V�?EH�>��=$׀=[U��,�>�fk?��<J�=�Y?�(�>���>DƲ>z�M?�,.?B�?��鼬�ýXM�� ���������j�=���>�>\>e��>�#��W?F���
	�c�4>�@ǽ�䵾�q>���>_��>0�\4�>��:��*�B��>~�?S�����>��>*��>�����>jC��j�����n��=�F<\���Ym>��>8��>-�?g���}<�>�%��Fp�>��t>��=�m�0�:?�?v�>���>w;�����>H���>�޽��W>��>�G?�S�>���>��j>J6�>�Oݾ�շ�Wo%���>�V�<%>�.=*aD�5����r>z�=�zh��`���N!?+��_u��¢=��ѽNPi?Ц�=�##����>�Q�>M�����v=�k?��=;��=�G�u%?���R��<'>F'7?��>���>i`/=Ka���S����L�>�UϽq�>�E�>`l�=������������ț��o�;-l����>Ò����о��!�����{�>���"��5V�=�⍾ġ	�I>˲?@��>S��O��E����ǽ
��<�7>��=ވv�1!0>A/�>��>�G=D��RP��׌���a��A�Y�7��n ����<��Y�ۃ�>�(l�L�>�gԾ����|�c�C.~�:I����=.�>��I�%�p���s>���*�>��A>Z�/?����_޾/R����~�>iG=��g龊��=�Y�p���*Y���龩����X�>Y�H�n��>Ħ�9�a޽^������j�E����w�p�?�yn>��?�W��]>m�>�:�>m�>N��>�K˽�B�>���>l&��p˼�������h?ymF>����d��B��٘&�K��F�>L�����>��n��?܉�>N�'��J?c>򏓾�����+^���=6���>i}������2w<�]P��H�`U?1�>���?GD>�>��p쨽�%�(׿�Dv|>T煽y�?�����>���?�þ�p�>���>i�=�;��&G?z�,�>����@g>�m�&"�3?l>k�	?��2?����4�>Z��=�ջ>����%=\B�>>�{?��>:R+?��T��0�>�==?���-�o�����[>&E�=g]?��d��^�>��.>���?����$���p�m�?㾷�7<��w㾄�d� "��Z޳��*��g��>zx�>A�/��\8<|�;>?��ʬ
�Շ�4}��5
��Z�=�W>�)���f����r<���9/���������۾����*C=�8>� ?�>���>Hz	=W�q�i��A�z�˹?+��>���>?:��ӡ`?�>Wd�>�>��>} ?�-v?�h�q����,?���>��ɽWf�rQ�?A}?X;��^�>E�I=��>��)��X\���X>#G�>�3G�7�ӾoE���'� ?0M>M�/?���>����C?��>j�Ld8>���>^Q�>�?A��>���>�q?�c	>�]�=dQ�=���=�k>>@ľ��>�t?p/Ծo3�_���Ħ�D=��?����>,�<?
�>���<Z/�;���?�R�>[z콱`!?��>\?������>ӥ0?w>ͷT��g=ޗ�i�U>�B��|՞=q����%���&����ܾ!zV�̸x�餩>FPl�iaȾn��>���>U��ry���
�j�>Ab�>��?���i�>�蒾� L>X-��i�þڨM���=��u���AϾ��57��̆>|���6B,?l<�cp	=�V<��>���<YF�'@�:�7?���93���~>������?<�u��������g?�-5�3���?Γ>!��>=�r����������?���GH�����۾�?[I?_�\>4�~�A�?�҈>�X�=�"�5��>I��>bjw?�E��jA���5��C2��r�;�oA>㡾U?=1���傾	ʼ��*�p*�����-���z�>\F��}��>��t���^?7��=�S�>3i�%m
�=v޾�=�aM��+4��(�>���*���﷖��,f�ܚ6?�f�=M�ȾgY���b�>:J?wXm�kRR��8?�k ��y;���=�l�>���>��>L�j ��<��#��>�⋾�eU��!3?E�>�[澶���8�h>����>�o���۽�p���r���ѽT��>�Q��?	�>}�W^��9��;J?sE����ʽE\&���!>�g�y�����^�>�R���G�>ԁ^�N�>�͐�B�>���{�h��I�X�X� �E�=�p>�[?E�q=�4뾺��>Z
{�^�z>>G=?�m@?����Syf>�s?�5t?\�>��)=e��=�>��7�Γ��V���d*���B?��>�/�=y��	X�>��?>r.?��:��aK>��1��"l>�t���>�1��&�0�(͙�س{�Ń�%|�>���>�u�F��&&�?"=�>����v�>8+��:�|>ï
���/���M>��a>�����>C4?��<?�5���7?Jbm>�㊾F���~&,��h�>T>y�A�f>*FM�+H�.[нZ��=˦s�4?�u���<X���T*=d��c6)���I��&?	M>2>�=Ͼ���>+��>��>���m�<�(<�=lU=�8`ž
�=&�;�����?:�?Fa?�F�7la>q>B=>yL�>Z�'>�x>��u����X���?�J�����-R��@ӓ��>�)�MJ�>���=43�>�Ї><ݎ=�>X�?�i?�O	:c�?��u�i��^�C�9�����Ž�Q�w�4�1mV���B?wm,?�z���-�=ĸ*?���>&F ��9�>kf<+=1�� .=��=x��ō6��Z?+1�>��>:�W>f	?x��?dd�=��?�
>&F<H
J��n����>�BJ�h@%��콱�d>^{7?�
�>4:p��즽K�?t�]>, ��4��>�}�>�0�>�k;Aj7?�D ?V��=�� >`�l�d>=�� >��潶�>>��[>�*M<md�>{�5?��[�%�>����߻=v�`��*?=$K�����;�ц����#>���b V�,V�=__������4�7��?ʇ��V>+�z��">��y.�żþ����9?�k�"wp?ֹG�����>���>���u��̊�%�?���>��>���=���=Ot�e=�>�[q�2v?�*(��j^>��
>P�/?s/�W��>��=R|>+F��±��*4�Md9>��Ļw���+`Z>��?~?1о�K�>V=?����B�E���W�����r>q��=m�)�|�2�;X���=�7T��l��k�G����h������	���>� �*�~^�����=���N��XK*��@���>[���P�����X>9���q(��$���=?�:@=�0�fEB�A! =ء�>i_�>��C?��S�إ>�(���&>,f���z?>"��>kq?)��>�9.?����P3��]��=<@�>^e��:M�@�w>7r?�c��컦�@!M�Z�Ѿs����L��}�>#>c�>����=��k>��>��9��d=i��<6�1>z�+C>b�S?�u�Vo潦W���/=t���AN��.z<�Z�>���=C�ƾ��8�U9?d�+?����	�ñ�>�ƹ� 	����/��*u>Ǳ$��Br��ꁽ�y�>����V0���y�g�Ra�>/T�x#�M�?��o���,�7��3hL>��>f1������9f��=ɽ�7.��=����>.� >�>����{w��
v�>N��<�zD�r0�>*󽷨s?�	?������d
K>�\���"о��J0>T#�=�Jս�xi� w�����=j���#����3��(���-�>}�K>��N��>T2h�e��G�>�Q ���>W�Ӽ��.���y
?�����?uB�<��<j�=�=?���>៭>��&��m�>`ճ�L�l>�v>�cy?���>��|>���>͞?nn>�w��z�>�$�>G�|?�jq�O	>����/����&?�b?�QֻQ�=�����
3��kܽ�����Q?�ţ>�}>,�<H(̼�BC�7��;��?l��Q��=�F�=]?�qy�g�K?G��>��>��>w{Q?�i���@�>|=�	�=Y_�>�+#��p>�.=J_���u���>'�S�p��/L+?r�h>Z�?>I;��ɼ����>���>�(��kB��mӛ>L�S?�F�>jJP�t?j�>I�Ͼ��>��>tu(���y=�>���=z�����=_$?���>��=�<ֿ.��Iܯ��X���-�>����*�U�I�����?��.�Mо�g�N<�$?bh��(�o���!2�?�?��?4�>K3?~�>�;���DE�p-S?�0-��s
����>q�>���������>�d>���b�6>s�"=~��C#��]�u~Ѿ�k��B��>�m5��>Ğ��g��?t倿�ɾ��"�B�� ��d�׾d�p�ۺʾڂ����=�>�S��X>�#�����>���?�=QW��H��?q'F��E�>cf���X���>���7?�R]�b������=��>eZ��{�G����?��J=#�^�9e��P1=��$�s]پɻ$>����B�_&!?�������J9�̵�>CC.�#���l�z=�ʪ�`t?�T�kN!?�)tn?�B}>p��>��,?�9�?i��>��#>�E<����e����J��Zj=4�h��u�V����>+��V���Ȁ>a��>.�f=����#�?\���f�p���9!�>s*�?x�{�l*�>�~��O�̾?�<?�x*�_;V?���)<�a�|��#�9��~ǔ=�Ą>�h�h>�� �ps,?�A?�j�� ���?$>��?�2>���&Z�F鱾bw ?���>
1h>��`��LS>�Y>���=17�+r��-��J�3F���\�>8.վ�B��x}3�Y&-��6ξ\���f7�����n���������gJA��Xb�o�N>��>xkR>�e�>�X���?�>��=��վ.F>
WZ>$&S���y=��Ľ�9�>rD��˦����(��fy>�\�>��ܾ)E
�E:�>*0?5��=Ep�>�:'?Wd2>[��a��˕F���:5e*>4�>%�=�f��Ъ>k�=�>5?dk�=3᧾�'�>9��>�N>_���������>�k�	��4?Fξ����H?]�V?����j��G�DP?y�O�m���CW�=��>M�,��.��#�>�љ�r���.��=O�ѽ̪l���.�K��>,GF?O�=�)8?C�]>:�J���Y��������81?R�v�b���5'�� ��>�*.?��R?el�Ԋ�>Q	�>�O�>�HA>~m�>���?)�,���>>�0�>�O(=Ƞ2�������<�����>Y οH6?��J���mƿ
��>+� ����>��?�I���<�>�羫@R?��'>��w??k=Xg���?+�U�l�n�§��rs.>��t?�{�=�;�>)�����%?u���eYN?�Yڽ��>Dv��#YS?�l���6>���2�>4�?x���� �=b��?�W�>�mh>n��g/?(��>v<a?dw����@�<>��>6�+�E�=+p��p?o)��SK��༾eSY>7�h>�L�K�����ߓ?����Ƈ�=�1��S�����@�-�>t=�>r�*?�(?M->��ӽ�x?
 �?�:�=дP��ܟ�������h�s��CV#��ﺾN�\�G���%ì>��2?R��= e���>W!�>����(�F� ξ��>� ���2����>D�)�$�=�7>;𷾋� ���=uv�=����ڻ�_�v=���>�O�3�潡�:a�<�a��Es=�璿�<���>�d���U�����O1.>�7_=�/�>��L>�!4>�
�>�{�=~�f=�e���澗����ڤ��}>�J�>{�M���ƾ�?�>��><�����/�NѾ]j��"����㾦0>g&�f��>[�.���<�&�>�X����B>YꋾՆ��%�-��	�<��>��$羴�?~�<K�?|�������4?�0��SlٽȾ9>M�>�M�h��Oǽ�^�>)�H���>��>+�S��?��?>�^�r�P�&�C=2�S�s8�>1R>i3��(�G����M��|2������v>� ����>ࢶ>����5,�����??�@�o.��t �9A>&*�>A� ��u>��x>��>�_��s��>��߽�0��%E>��	?@Խ�8½i��=nҽ�'g?j��N�?�~���>g�>�̟=\��>�3��A>��=9�?JgY����>�aüL�?��������ZL����
��>�	�=�g�-Q/?��?�>�Z�:Ѥ=I(?��?�݁>�Y���%� V �8Ǽ	��=X��>B�>����8�/�8.?�F?���=O���>��#=&>*پ���?���=ٽ�>y"޾�R?����C?�D���]�>���H�?�ɾٓk>��=[	?�Y�{!���$?�2G?}�n>�蝾?��Q^?��W>@�� �����?{��=��*����Ig�=,�?����@�>5N|=�?N?Q쑽+�m>��&�<o���*��?&�>	�,�5b ��0当BG��A ?�v?� >?V�e>\f ?#����c?��o?��oD����>%�4��2�>��>�����$�\i6?h��=g�м�no>,ë=u~��ٚ>�(a����>��>��7�EU�>�(��1}?e"�����Bƞ��>)���XB�L$&>.�?髊?Őo< ��)I]>��2> �.~�� ��_�="f �@
ľ,' ?lhm�5�y�a,�>:�?��;(?��W�ս�Ͼ��Y���&?c��=�$�>hK:=WY�=�����/���>����[��>�q$>d�>�M���l�=�6�?���>�0>������=?;�G>B~?�n2�ʍ@�=�>���>{�)�]P�=D��4 =���F�R�=�?�>������<\!?U��>����p�F��gD?�ܾb	��)v�>����3[� ��>J����SA���}�w >��-=zDξdK��m�4��Pe?�r���.>&륾N|/��t���e���
>�����_�>gL�rV��	�>��7����=-wJ=T����k>�h ������&�=��N>�ԍ�rgO�}�E>�'?q��>
��n�9>�v>(�h>CN�=+.���K9?���@$�2ݸ���>4�0Yn=�y��}�>��>�6��]u���o�>�e>�ܯ=�?`�k�?yC?y�~>b?D�]���	����>�(9�+���ptl�������>��[��н-��r'?�U��_Ƚs,���
?D���nX�F��>!�M�'�H�ז
���>� E�͔��̕���
�-p�?��࿿�x>���.���b�>%�� ���G���o�� ���'h@�j\���:l>��'?�Du��H�>{4?n>?oA��x��I���>Ù�>���8*�}n=�[S>7_W�B���3 �<��Y>'����G>��#>D_�>u����>�I�=��=�G�A�S��o�>xW�>�_�>�\��t�9C?z�*���B=�p�-k��7�?L�>x�>�>��{�B-�'�v�|�?I?��4��ˊ=�B^�~z�� �޽4���/]�=Ͼ��]��iZ=dt�=���8��W�(��=�lA��}"���/�(F?�����6>�Ga;�쾾4	#>3!���\>j�=��5ľ��վ�~$��??�tܽ D?g�־T����e?q��>����	�>�p&�^q2?v��� J����
|?R���r�����G��O��j���tw��\�>7����/��`�<�̃������֣�;H�#$�=����^=�<���=0I������ͽFCf;�*ѽbă�v��<��=�=>r�<�^=6>�=y;�=�B���=K{�=Ҋ=KȞ��>p�<�i�=1Z��>�Җ<v��=� ��V7�=Q��=w;B���!��->F=�E�<g�ڽf��6�����m2�=���=�[�)s�ș0�]�-�'��<xD\�+��<�i�<U�@��RE�߱�=��[�A5R=oV=�F�ޢ5�z@�<k�=Q0սp����c��=������PV�=�Do=�
Z<V:�:��=o��=e{W=�s�=	j�=�U�=h�9=�d�<GI=���=�m��Bq<�tB<V��=������{�=6�>�Wp<z�<`%P��U��e��٭9="�=S�����.<�WO=���=�=������F�D�3=���v��=f�\��.��oO�`@�=�R$;4��2p�w�=��o<�><������=����<�-��;��=��<�;��-~���\=���� �������x=�M1=O~��x���=���:���� ��I���(��:$̽U���\ֻ�X �x��<4k���0B=5&�,���ҽ���q�f�:�3���B����f=��������8����=���W�<=���	>;����Ľ�5���<H�Z���R=�=��c���X=g�C�r��<>7��Ww=�j�=J���z =���FǓ=j���Ný��]=�ӽU[��=�����ở���=�#1;�o��%���r<�!�:���5<m|<��k���Y=)Ը=� )=7)��,�<�Ǽ?�=�ȼ�Ŭ<�x��Ɏ�]�==�����{���G="��='Z|��p�=�G�=ok�<-N�h�=�9)=��b�E���s6���<�<N��N��<�p�<���L�w<>��=��=Qf_��V�<d�;�=��Qл.�<F����<��H�g�
=��� �O��-�0�&�>!��%��^�V<��G>��ǽ�a�=�.�U��=�*����g=G�[=g��=����ޖ�={ڋ�a��=������0�mB�7^�[�����&���<&�W=�û�x��<:>���4E;aK���=T�x=�h-<���<q�۽��v�?�=<�\�=�2Ѽ��l����=�4=�^�<�S��V8�ؠ�\�{�_��0�~��Ճ��8�<q�S=_\��Q��	ڽ��>�ۆ���S��:�� >E����=ɀ�={>l�<��D=�W|�p����<�=F�6=���h�M��i��֣�<F�<�Z����I��p\=��=d�н�V�&���]*�*�ļ�6K��&���	<����7�<^�Z<�Q꼙�z�-	�%�L�6�	���[=�&�=�1z���=c�ؼ��i�i�@�|l~=.pS<�)L:�‽��L=M�=c�E=i�;3�#>�2�;8w�<z����,��0�~�^�;�U�=�|=����Pw�<h��=��R=��z�~��=��N=�
�<v]P<�f�����<��=�٣���=�P�;�2A=tA��/^�=|tk=�(=�.����=�&=pȮ=��`�u�m<��̻�!�=H̽>b=:R��ʠ=�w��A����<Cq��Oց;�Ř=U��=���=f푼Ô!=�{=�g�=�(d��[�u�\��˳=��yZ�<��?=c��=Z��=G=:w�=��=5�g=a�h��r�=o���-=���=���=mh<-���zJ�=�t+=�:�X@=Y%R<ܚ;=���=}�8<�u=U��I��=�N����<�e��"=Wa���D���>���<����b�6�f`=��=��=��E4��6=l�=�^�=��߽�	=	��=������<�W���׽>n�<���"��հ�����=\5=B��<�~��r��<͟-;[tc=(F��3-�M.�%	o=����|�Ӽh�Q<G0<��=*~�=,=�;�轾�J:��ȼa���v�$�]�w=��#=:��<B�����=�a�=ƭ���:����H��b��\(7=U;ǻl�"�4ǖ<8�>��<��;s�H<�cO���4<�!	�V�I<	� �~0<P��H/�yݼ���<������#�l=�`�4~���c������N<��&�۽�{;���x'�ɏ��ۭ��(��;հ��9��<a�<v��=����6��ۊ����;�z���ǽ��<K���7<�}Y����=���	s�-��)Ǹ<�u;qQ�����}�=�*��2O��X��v{��XQ�G�8��#��K�}<s�̼�&;I_�<�' �0@�;�k�'��������e��V��!�^���S=���=<c�=#�=r�*���>��޼��=�ܢ��������6=ɠ(=�n;In���=Ń�=�B=�H$�O���/��=�,
�+�������D;pzA<O�ʽLP���!���c�X��<���<�<��h��=�Tx=���=x����=)A�=S �=W�x��-��o�=�&=�."��(�G�@;����M=ks=�{=�+��1�=a�=$w���`z��4=�=��ü�1�m�#;Z#��t�Z�/�ν��6�M�=�Y�<LB#>j����N=��n<���=�$��7�=�>��=}����k =�R�=!8=Ȭ<zG��þѻ!i��E:2<���eA<��=��{�\�<Dg�=���=�ه��-K<�%=�'x=-N	=u�����<k	�=�]��
�~�Jt$���=�?s��ú�E�+<#�=	��I��=7|˽�|=G&|=|8ڽoݏ�����%�����}|��V�<�-���-�jΛ�)��u��=��M=��=,�=���<�ʘ=��=��=��<'�<�{�=,V��SPE=��=��S=(�=�l�=$�<iR���2�0�=-�=I�	��,��ϧ=��<R:.��1Y��MI<o�4=�d!=:��磻/����ڽ���ɺ���=-��=s�>�ve��m4=�>�F���_��L�=���=�ZE��F�=�vF=���=SV����*<�����d�=v�:<p[�=K�R=.��XMA�Qb=�'==��[=c��)WV���7=�@ǽ�����<U��<��t=��X��E�=��I=�S�=���<V��9>=[=��ü��="�=�t=�Kҽ���d鑼R�Q���j�ZjI=�=��{=�*l��e���=�=���7��{��r��@��==�D�<�$�K󵽌~�<�>��=2�cw
�q��;�u��H�����hM�<�r��A��G�?�-��07=C��Խ��Z;zƄ�ӭ�=ﾝ�Q�=E�+��X?=�O��KQQ�h��< ෼��#����s��<���<e.V�US��4�Z<"�i<���=;�=�ǰ��Ke=�����<&zk<CTE=*Jw�O�6���.=��s=��=B������<��=��!>N����ֿ<��>'Y�=8[����%��B �s�=���:ȫc��ef�'�x�ѽ��2�o�M�e�ޜڽI�k<��;�H�a�\�R��<3�cr����D����9�U�:��<�Q���N=��<�d��X���Eg�<��+�
��m��,t<=���E}E��n��{���{��?C�=�"�=��;�:�����<��=��Y�$��1'=GO=�i�����;��%���>kZz;¯~<'_�ioJ�Hz=�*���h��1d.�;��=eŨ�� ��p��@��<&�<=�Q�����?�=Z
<�=�%!>n}�=e�J=��;��;�!H=�7<����V�<�>J�;���VZ}���=�%>�O =p����*�=�IO���k<o�^�ðH=Ѣ;D
��Tx~��*��ʠ��K����GJ�;E�ϼ`Ľ:���=�q��)������h��=�$0�����"����e��ә�hN���*D�~>Ժ��/���H���TU)=,=k�;�ǒ����=lC=l㌽1ꍽ�P�<�p�=O6L��mz;�<�<\�=ݣ=��"���󼼇b<^�B���'��=u��s�=ef�=�f"�Xa��*��>�=�@�>�������a�FJ9>�	�E:/�{�=-��=���>��y��%�=�4�>g.�kԾy�5��ޡ�=M�d���>�1h>gL�=�b�=�f�=��
=aJR��	`�vS�<�T,�C�>$���]q>�(�\��>i����3���3��9�m�p>�=�=�͊<��3?��G=ZI�=���J���,�����1�>uH`��7�=o�>"�>>l�Ⱦ� D�Ƞ�=`���-�=X ��=�a>�w�>[Ͼ?���v<�d����Z�<[�<�;>�'��F��;�
N>0��>:��=�:ڻ��ϳ]>r����j�!�L���=� �>dx$>c�I>&>b=W�I� �|\=�撾pR�=�l�$�??��>Z�{�]�彁������@�=��Mо�ɾ�ļ�D����=.��>��>~^Q>S�I����~O��n[��/����ZN�,Bо�"��@��c�>�.����L�I�*��=b�3>��V��3��B��>CB�����=P�?��Շ>T����]��Tۼ�˛>H�����I#	�$�=�2�<Nɾ�6�h�-?2nӼ_>�vt�T^=JK>��>�e��p�
��Ə����}K��s���+>b�]=��8����=E�t�tT��x����s>�.�W�7�Y�A��b�>Q_�R����`�^>�>⭗��I�����>q)ʾ�`\�~G������$�>MF��M�0�o�"�p�����>�F�=�8�>p�O>:S0>�3D�QG5�j9��������V8�>񜈽�v=lS>��b>Rl���p�G�->d��6��=�>{�&zl>�i>�I�����=�?�>�\b>dc{>��t>h&��y*�v~+�����}�������콽��>#~?�����C>9���=>���=q��>O��>98 ��O��Q<m_=��i)�N�p���U>���>"+�>�h>�d>����ҭ�=T���x���뾯�e�\'=r�l>�ŕ>m�F>�1=������<e����Pd`��e>�����\>��a�>O>���>�$Y>��=z;��kJ�>��b=��g��>�2Ӽ��M>��"#=�m�����Ħ�-)�=Ϙ�>���>��>�	L�6�=�H;����)��<����;�>�=3s;=ڱ���hx��щ�3;ͽq֘���>�5=�8	>!D޾ˍ�@�|�u�������G�=�M�=C�?���=������=�iI>�
���������Y)�>��>��>Cp=o;�>ݽ��=Ӝ��˧ؾg�;��<Vm�m��e����@>B	�=a|ѽ�	8�`64���=�M��y3���!>_�;:�P��xD�!$r>�}[>]X���W>�I����=ل|����)ϳ;���=��ӽ�o=�-����=���>LS�>�]����^�=�v��2y4��sd��i>U��>ֆ�>�g/>�;]>g���`Ͼ4Ǿ�a�;�.>��>hP�=�S�P	>�S=�ʥ��M�������I>u�/<\�'>�����P>#[:>�nJ>º���pZ>gP�=�1�=����Lپ�p�>�F�=�4�ׂ�>c�=9,�>������ɽ�;���wC<�eQ>�ʱ>��>#��=Q�>��>����~����?�!>�	?r��=�d>�-U=w�w��W�Ou<�"�>Xs�>H�?�~�=\��o��=�ܾt �\Ϳ�i��=U���>�l>p\�={�=����h5�>F~
>�X�ޔ�������K>���H����ׄ>�F>�e�=k�Y>}kS��w��&����>i���}5ؽ^<�=W�3=�um>�,�J"�='{7>]j�t���`�<6ܻ=�հ�� Ľ����%��@�<��D��W�e��>��=8Y�=��ľe�ؼ:�g���,�L��Ë���P <��w�$e	�����uyS>FA>קZ�?�=G�<�O{>�ݺ_���%>"w0>?��<�T��2Z�=�^�>pڵ>�vq<	�M=ms����X=�+��!r��^ �<�*>[��|q;>�|
>�;?
~�
Wݾq#��IMe�ۡb=ﭼ<�Rz=�m��%�?f�=���˻Q�>���h�=jY�<���=�����
��M�("���&��f>�b�=�z)��=Q�d�@��>wԾ>���=[>��=M�=�p�>��ؽr�>|���I ��Ad��ؼ�� ��ў��.#>�o���h=���>�־&�+/�OPI>��+��u�<�� ��dv>��ѽ^���I�g��U'�YV�>&���G�����h?��K�f��=>���5�<���= i��}(������,3W>A�>賱>��>>kU��/c��e�����
����{�>̮�=�L�>���>ǁQ>��6��]�=4�<�P��'�&�ۖ��I�>V�>�>7Cb=�H�>�Y�>ժ���H�=��>�@^>����t�O<>U���:�==zn���>u>-܅��g�������ĵ�"�>z=.>{X=g��K�y��=�j>�8Ҿ�P�/G>q>!=��/�����ǁ����==L<!԰����Y�ֺ�B޼�v�Y�����>��=	vx=��n��Z���ޡ�I������f�o��>�N�=ϫ">�����%�=Yt9>��=��&�L�Sq>e2�=� !�gjF>���;jV�>��b�j�>��
�-G�@뾁Bb�)��>\%�>iq>GӋ>��L<,�!�U�?����1��ួD#>6�o�
">$�>���=#1��z��>R�=��%��Q���>] y=�^>�y��9�>�-3>󎘾"�v=�7�>t���{�u=�����L>
��\����D�,_e>�ey>�jh>�{>���>�4�=��=PV5>�E>;h">���mŽ�Β��>�S�>�"���U>;�<?�%��sK>���9G@>u���B-;J�6��?��"������Q ��c"��d>5�A�ԓK�Z�>P
Ͼ���>�3�����=��>��D>7���6v	=��\>@;�>W���)����=#O�>����y4�<�l��C��>�&��K�>���e���;��ed&�P,�>���:�q<D�>��=A�c��Up=1��ٗQ�!����ɤ���i>�б=�}�=s j�#��>��=�n4���T�������%>�#ü�5A���>l;>b��=����8F<UEs�&lǾ����?>�l�=4U3<M�}>��2��.�>1qy�������=pB�=1oU��E�>;���n��*�����b>�n������<���<Ǆ>��#����=C�>�q��[}z��*���ѾQ���|�P���q���%���>��=XK;U�8>+�*�r�>�Vž�����>��;�ju�><���"��=�,Y��pL��)۽�>�g >�I{�+�=?�5�y�>M���7� �돂>C��>U�e��nY�{û>F{�=Yd�<�"��a&�=˚E>[��<N6���P� b5>���<J]��3Ӛ<f.�=B�4<V�>�|d��x����½���>:�8����+O<��*=��>=�+��i=��>׭��,�����c�>Z�Og��^�U�^>��i�DM�=P��=!Z�>N�3���=To�>�I����6���v��0������=�}>=�X=)��=�	A>ܴ7>7Q���]����<��q>j�Ž#��>��'>	�?��f>tw����ٽ���<>��]��ZI�yG��Ⱗ=<��=�`����<��>��4��ʁ���X=��>�4�>!��>a�>m�>m���8�[l�ET��ߤ�>�����W�>�h?�n�о>�����>*!�=A�ټǽ�Ώg>�ʽ�����P8�&нJ0i>c~*���ƽ>I@?H���%��=�W�-|k>��G��ܽ$zo���Z>�+5��`���JN=�9�>�JI�񫩽��9?�����$N���� ������V�c����&�=��=C�-���$�r�:?�{�<�%���.�Qje�}�d>|���<<唸=��^>���=��@>�G۽#�l��+>ru�=�{���y:��`T=��>�H��y��qE�=\�>G�?���;lF��Q&=,o>�[�Lw��J}=�~g>� >mpd��G"��R>\�u�l^R�ʽJ��B'1>~�>��Y=l��=4v=Y��yu>y�;�����>a�ا>����졷>���=��ľ޿ܽ;>Gј>:JV��(^��ޑ���> e��uy=Ʊ�>Ǧ�>��t�V��"1)��Ͽ��ْ��%e>�2=Zf	�F�=��E=���Xħ��0O>S��yU�=�s+<tY�<栂>!��B�<�:<��e�q�9=Pu�=�̅>Ubܾ�5X�p�⽥�>{�=7�jd�;�	?�;��?2��w�=s%?1��=�`>��<Y~�>v���g���<��>�>Ȅ���P���I`��(�=�0>�ٽ���=��n���B����=\9�>}����E'�(O=��?��e����=m|�>��>B?��oƎ���羝�Q),���>1\�a�Ѿ�f߽�7?Y�,��!��B����>�\|>eIK�x��ɦ>�>#_�������?R��.ʾ�����h?���|���P%���gQ>[�>���2$0��n�>aɎ=h�p�����!��g��+�=J���_��=-p==�>}�轝$&�I�K���@>F��-�=�5[�����`��<��	?6�X�J�����߼��>��/�g辪��;HH�>(Y�>9��������)>�@#�D`4�d*�4ޱ��:B>;>��+���b�!P���g>�f��d�=�W=7��=����k��! ���
i�0�[�� _>Q�ܽ��ֽ�Z�=�d�=�j����ھ�lB>�u�=o՟=і����;>�f>1�W�8��<.�=�f�"e3>���=��>@�5������8���v>�GC��2����=Ϧ�=�*�>'���"�r=�0>lS�>�;�]u��K��>��2>�֜�� ��>ZPѽZY���!S���>�"�>���>Z�>$K>2,>�1�=-?;8���ɵ��aQ���k>�͎����>
/�>��y�����G�5��G���,����:�>��<=��i=�@#����=G	�>0Ӳ=$Ɉ��1F���d>4��>8�?�>C�>�h3>�<��+>�_�;��7=�����q���[l=f�;>��<>��=��>��>C퓽:"�<E�>�B"?��=K����9Z�Ǿ� �>?��=��>l���0�>6�=�m�=�l��溼���-��;I���+.�s����=裰>)}Ⱦ��'��2J�m ?(ڥ��*��[=��#?��>D�4>
��>�#�>w��ƵF�B۽�h��H`=L�>̨>La���}N��]>�H>�����1 ��^���R�ܾ �����= �=�B�l`��OT>�t�>�J$��V=��%�FA>h����۾EG�q���Vj�>�$�0?���"�>��7>�����PGN>�f��P������멲>���>��?<��>W�f>�/��"��o(���F����!>�{_>�E=�ӭ�p�=Q�?=wj=����'����@>cQ�=��Ⱦ��m�>K�>�~�=�I��|>�1�>7�E=:@���̩�Jh�=�.>����?�=(ɂ>�g[>r�žpKn<���������>��#>�=��G>^��=��;;������>��ڽ�l�>`��=a��=�$�=�٩>��;E4�=	���������=��]>+J�>�/�=�V�=���=C�"��q����	��J�>Ĕ��A٠>է=>�Ƽ>���n��>���>1|������C2��J�=��.�#߂��}�=p�=�[����>�����m3��7�=;b!>���r9��?��=A(E>��>�,���H�=��l>�̰<*��;l��=U��>^��=�= �f�>aST=�N�>_"�>�ֺ=ZT���%��=��Ղ�C޾�|������\ѽ=�Э��Sk=�b>X��>�=y���4���$<�´=�c��,
�6�=�i^� ��o���ܽwI>p2�>��k�3='�4�3[�>�}��?�b�
��>(C�Y��=�0>M�>����9���M��a��D��>���=o��=�]���~�>[�4>.( �i�R��8˽��=fe+��3������A�x��==I��jBb=�5 >��u>?@~��W=-:�<m5�=�=��[A��p�=��"=`�'>���=�c�<��=�������m�����|�-oP���]��
><��3>�xO��c��t�v�:�?�;����=��B��0(??�H���r���~����=�KQ>��:�g ��2��>C��吥�VLz�O�ټ�T�=�5���Ӿ�����檽ŀ>�-;N>~dd>W�ɼ�Ğ�ş�[��EF�����+>�M�>�T��E�>���q������G�>ol���½!]���"�>0�l>�>I�>K	N>��@>~��H�0$M=�VZ=fg��V��3�D>��=z�=c�����=�"A>��y���{�=����b*�>,�?~*�=f1'���'�$>���h&����q��j)>�V��<������ǒ��+;>�i�>�(�=��;E6����>%ia�k�:>�1��p�>sL�=� ��M �v��;�X3�:!�K������>��!>L��=�B��Y>�?\D�=a����F�(kT>�6>`پ��=VA�>��><Aདྷ[(��bӼ�̆�񗳾��T�iƒ>� ��-x>6'�>��5=�]��Ӏ��.�Id�%nf=�׽=��_<��ɽ�?|A�����h�Ц�>D7.�V9��R}�i�>�.�="E>���>r�M>�>'�F�\�Ù�>�G��7ҏ;.�Ǿ��;�=}�j�d�K���L>���>nA�>|�?���>�۽�+ս�̼�(> P>�>�,ü�9T>Dgg��_����=��N�Y�>�/�;����F���>���=��=��̽���<c��BE�0���v�=p�{=���;����`�=�૾րp��������2M>�8 >�H>��[C��p^��>�w����r�h={2�>����v[���r>�`�>SlK��@l<K>�Ť�ig�4�紲>V���Z��=`�p>�rl>�7�r֝�����λ��tg���㝾��>#�>�����l��p�>���>=a����� �u�1>o#���s��I��=�7>�o���w��x�==�>�-���v�����=Y��>�^�Q_�=�����A�=��<�ݜ��D�½���"���ՠ>�#���;��o�<v�/>�DԾ��ξ2��=L0#>�^�=?����;��>k�y�@������BQ���@��=h�+��j�<�I�=�4>\�8��:>��5Q}�o�=���R�>T����=�0��|�D>B�ý2�'=�'>[v�>�H�e=�Gν۲8>�YO��n�u�>�n;(G���о���=�fJ> i�=S���p>�?5��<���:��p!n>pc�=	��r���h�=����Tg�>�E��>N6�kt=�/a>"&����AV�=��D>��(>C���B=�c�>2��y�	��!�=���>��8��[��<�H>"A���:����<��>�D>}�����G�>�);�3�j��;̽��q����=��H��e>��ξu"��������>1L޽�yG�m�2�P�>�p ���>z�>�0+>��>eL�x�������Ao> l�£,����<�3+>q �����P��x��>��3>N�< ��=���><.�=ii�=�<�>=�>Ҽ>��z��G>5wO����=P�=)И��>��:L�ܽO��8h$?�3�:�\�=i��5*/?k�{��y���f���=|�=;ږ��Ś��Ծ>��S�E��bH��?VҽC���A,ؽ:��>��P����M����>��>��S�C�b���>fg� ߾&%��+�x���<���\���p�>��<�X�=Ƭ�b$?�$ ?ѣ�D��ӻ"��8>m�ŽY��'�=1�	>�>�׈>�L���-=��!�Q�=����Վ�/�ż�]>��ž��e����>Y�2>�?zt��aU?v�ӽ-����ߐ�f�x�ԝ�G�?W�v�?��/U���Xl�>�����=&Ɂ?��ȾA!վs>�P��?�o>)��>K�ͽ�?U��(�*?f�>6E�?�ظ��!>�;2��=|�=? �?E�I>��>^��=��u>17ʽ���<���>�Y�=3|�=�b������O���TT=ko?��=�?�
��Չ�>�������!�>'�h>�Z�������?̾8(>���>5�>=��|Z?a�?K�?*��lW� j����>�x��k�Ͻ��v*f>�A��ڀ=%̌>�G?T��>��>�e9?r$�=M�����	�^��ڇ>vޠ=Y�.��Cd=0�!��Ȃ��B;>$W7>mxG>�\�C5?Z9?f���'D>�d�>j��>]z2������u�>����^
��H|����~��n@�=�`?׶`���A�2���:�?�Y�����hh�q�?�?>V���򾾺��=�H�>�/>Z��A�?��`��9?�?b6 >�`��ҧ�28=`�?z��T��y̢�1��=���.��>r6U>
�2�]�$>ܽ>4�;��	=��U=��Ⱦ�ɾC:l��.?Jy�>�� ?�P�<�����$��[��e�>?��#�d���L�=%��>F(��6g��*T��ue�>}h����.U��ӈ>]�j>۪�=��
=#��_(�>$�?a�,��>�K�=�>w5��mT���:K?���/>���N�`�v�,~=s��>��¾��}>G�>EK�>�}���̤>�!9>&�>��'�#(�=-�>�L"��A->�?��>(�>���+K?�>�)$�s2ʾ�)ƾ��Y�ﾠ-�MV�=��L�$���/�>�w����i>� =��%�����q?Onw>۷��E��v?��3>�!�>�i�<��>T�A>�r?��+>��e?f�S?�ь���8�U��YS�ؿV����=�2?=$�,���j�˿��d�_ﲾ�����������>��F="*�>�p뾬�>{�>M>9�����=یy=#>��=]�=��>���<������>���c����geQ�Il<��#?Om���*>��*��j+?��V����
G�>��d>[�a���=>�>��B�Ts�>��>��Z>Ϯ+�T1�=��=�"�몰�.��>|�M�n;���g�?�<k���+���S0?�Ì�:?����=m��>	#O=煽��U?�d�=l��IU�>��?#|K>BI6���@�=�x������>v��?����6���l���7>��>{ǟ�݋����>��>�^վ�W徜;'?�&";cʾ%���(?���>��"�7YU��L[?�W��P�>�4>�6��N���C;�6[m=���[/����>�t$>�LT���Ǿl�?�3O�e�m<��=$�;�b�>c��>%2C?I�m>C׽�Jq�I,��:���~5?�dP?��?�*�>g�?���>��K>�%�=�A�?=r�>�^>�%6<�ys��#?���>r2>�5�p=�Ed?��>E�����>@>��?c��;�������>	�j=�
b�W����W��X>��?�!�=�:=CP�>�w̾�O�?µ?=eV?)$t?�O_=��3�l�g=�7�>�ư?�e?a�>]�4�2Cl����;Q�>R�=��/=m�C�⏓=�R�>�3�3>�>݂��c�?�>ت�=��j��E? �v?ؕ>{'о�3,?���0Ԛ>^�̾�$q��F:=Ь��(?\�6��~�����;/?�*�� 	���/>�b�><4x��qG>�?�[#�>�}�>�E�>|��>b͚<iZ�>qߴ>.���&�=�U�>5�K���T����>p�9>0����׽�>4���� �bˋ=L���:�.�<��Ͻ2�>k?}G�>9s� �>�1�>�;�b�q>��5>p��`��C�f��6[��Ξ�P��F�>E�>��'��c�>p߻�C3\��⾪N>���>�p��г����	>W��;������ξ��=��1?qٓ���кj
N>9�>l� >/>���ݬ��4��<X�>����x+��y�5�1����2��>�?Vf{>W[þ@�� �d?���=� �>�;=����ܽ�#,����>Ǐ�>�=?���Z	Y�E@;?S�W�g��Q�?�S��f����7K��k��M)��V#?��?k5?�����W��,���?�Q����F�����O�?l�˽I�>X̾ �<�7��[��تŽsн9+�?�m�>�������o��uν��=2_>2�q=�����\�8���tоݔT>`d����>q1�W6�<���>�ū=q���&�<Sz>I���*��	�͆?�&�>���=rϊ=�]>�l?�z���>���=_J�> �}��[O=E�$><�^=%�(��Ǽ�i�/�I���=���>��<v��=��?���>>�?����F��1>���T�$�U�p��R�>��9>�d�9(<��ݡ����K��>��>_7�>������=d���t��H�<P�>M��?�b�ص����>��l����Fm_��&��R�N?���>��>�k��F�>��o?V�?�߾I$(?�����߬>7�T'����p>�l�=T�>6�v?7a>�wx�2�/�ӞT���;�᧏>G�>ܱ�<Jн�n��6����	�V�>�������=1�*�:�6=��>�1���N�r�C>G�>���>>����X��:?>�bd>dU?�K�`?_�=˝X>ʚ���-�NBQ=H.�����@<*��=Ž�>�����Q<��$<P�'�^�?W�`>�';>W�)?����`�>�X��+>�֑?]�>2�=O��B�?�lW=�B	?�4�(%>�?�=��>���qj(?�??;-?����7�䰇���=�4�Ӂ>H�b���w���X�2Mj�����}@��FG;��?Ľ>?찹>�7��P�H��P�=�o�>��T�<��ӽ��|>k��!L９>��>�(�>��?���?
=�>,����T=e�)����=_$?1��<z��=�-�@�QB�-_׾6;ڽ�� {�?y�=�>r0T�܃T?��r?d�>*f����?c^���>7�⾡��}-%�u!�q�9=�>p^p=��ɾ�4b=q�?���>n������	��>^a>#�!=�
�=@~�u�����K?����dT����4Ą?Rԋ�:�|�k��<3>=(B�F��<Z�Ͼj��6�=����l=-��%|��`��F'�:hH�)#\>$;�=O��T�Ҿ<�?��>��?"�>L:<���=ξ���=���=�<��X�+�' ���.?9�?�<꽑�=]�}>�P#>�,g�ilF�^��<ơ���*�Ez쾒B?��&����9J�����?r�?h;�L�����>s��>W�>du�L����V��=���>z�ǿ����<h����?`��t��W���=�V2��e>,����m�>!��=)��Ad[=��?�O_��p��z�����>	�U�f�c��XX�=\�"�b��9��S~�z�>�)���r=��	?ȿV�,J���5M?|�2�;�=��L>�?� B�yR	�OD�V	=��#����>��>{Hr>�?��p�s�A>S�5=� ?�W�c�Z���/=�H�>����	����Y����>�����?��>���>�a����>_L>/�$����= �����T	<l�(�T�>�4H�ۚ�=֟>�?�LȽ�z�>"�΍�=T��x��>2@�=k��|��-��>�2���L>�1�����"q���
�Ҩʼx4L?lcM���Z����=~C�? �}�o���v��\ 7?b�=�-a�=�!�J�׽��<�a�<��)�bB0��l��������;��?���=��{S �Z��֌8?�B�<�ڽ�N�>�_ѽ��p>)�=�I>~�w=t�>��<�>��ZB;?���>{W]�ځb�7�|>�I�=�'Ƚ/��Zݔ>�<��s�K>geI�,nQ?C*+��}C>6��?f�ǿ�$>��@;Nm���C&���C��Gl�볠>3>��T��#����=6!l?8#Ҿ!6?��.�;��>
Mz>98?�3�?jBa�� ?{�>�#�?�X�7�=,?��}?��?x���3�:=d<p)6>��?P�>	'r>�RT?
yH>ia�=]Z]��x;�Z'*�䒣�2C����>s(��b�?.��?r�����>�?�>>z�=C
S��b�j;v>�06?�g:��8A���D�4>Z!?��>��q>u"��u�>���>c|�>y��R��Γ6>*?� ��peH��9��KX�k��=�/P?FLY=��*?�y?D��o:?Ż8?";�>���$�>)*?�Oq>d��ߠ��|�>_��>I�=��L��CL�����Z�>e�>\����=��5?eI>���d�Ӿ�t��ЧC�����亾��6=�d���`�>,��>�����+��鷴�GP�;�����⾭9���.?�'?�ژ��,�>��==8���ѽ�O���V�>v���N�YmR�B��I�P�V��/Ԭ�L�^?��5<���:NǾ��b>�M%��i� ����� �����D�>�O�!>���>�]I=V۾~W�ۯ�>P��¦U��+�H"�>/!����>�>H ���`�92v<(�)���������
V	���Z?oY��5�1��m�BI�>�/��K3Z;�1���);��{�>Կ>�6�>`h�?:���x,��3* ?m�;�`d޾���CZݾI �=��?||��]�P?
�?2�b��9�>l��>��>α��L@l���>��>xɾ)Fy�q�e>g��>�?x��zB?�7�>��y�6_>���NA��+�eC��ܘ�>"%z�ߡо9�ľ��?�b���F����?PD?cA=+)�<:��=}��>g/b=@Q��:�=�þ릙>ژ�>���>���>JX�{~9=��>ܽ��B�??Y3>�nJ�E�$͂�1���nk����뽟P?��A�y����y�a�=n^i�C�>�;G&����f?�{_=�E@>μH�?s�>��?^�!�b���k�>�����>o��ެ?й��+����" ?{.=��>�q;t>(=N>ś����H������>$20>X22�5R�>�FY�p�=i������5>U>�j��&=<3�W=�o2?���ؿ�>�>�>Zd>QW>�a��Ϸ>'g�s��>v�;=%���=�-�=r��}آ�/�T=0��E��>üK���ﾾ8?V�=�FĽ����'�9��8�Z(^��(���;�;���|?7�MZ������,>S>F���$<����� �>��#׺�/�?$�A>�\�L�@>��?<#�>WO�>�v�A�)j+>�8�N�R�ߌ>��=�>5�+?��>w�>bӡ���=I#	>�"��*>	��4��>M߷>�?��>?o�����nVɾA	�8)�ё�>����Sg>�F�?��=�8�Z>1�%�-F?8�'?v;�?1y�=��#��c��h�J?�{�A8��;�m?�s�=�z�=���> �,?�T>��v?N�l�1ސ?�>?���>4�C>��7�' Z�L���r�J?�L�Sj�f?��>��T>����u�e?��?��;?�\_=:�?
�
���P?n�l=����Y?8{=�|�>���>��	���?�A>����T��Q2�\�࿧^��X����g#?��'��߽f�?, �<�=륐��??l�? b?.�X��~?�w?/��\���?h:����:>uY�>D����p=��>\���j�޾|򋻙��>�R���\��:��=��$>���>�Z�پ��P=��>˘�>	޽X:?��I?TU=H�u�Ta'�\����.���P]�-���u��"� �R9��5H�� ?q����)����B+?"�潧�3��k���9?M�?�����=��Ծs\V�9��<]yپ�7ѽi��=&( ?�G�������>��>�$��r����?g�?�A���8q�<�x��xR��$$� �����W�>��(>��>��S������O>��>�q5<}7<�|��̽+�a�=�`/��Q{�W?j���}����=�"?�������G��C?ֶ[?����>Y>)V��ɵ=��?7���[����5<��X�Ⱦ��s������b�]�ǾuX�>/.>��=kE̾B�7���?L�O�n���}*��)�w>�YԾP���Pž,�?W�=c^(����>�#;�=����*>>�c��"�>�E�>Fl������V�>h���4�m����)�����=��#���2�>����n�>h�?4���Q�=?Ջ>�w?�3�;�9�+��=��>9��8s�Zh>���>J�b=7 W?��q���=?�~�?lMd���=�{�>4>#����/��>ǫ�>0JP�
E3�`�ӽ� �?�Yw>��<o�߾��!�¤L=~w�>�	>�/��?μa>X���c�*���+��������!?�A >��%>ϭ�U���f>a�D��S�>�u�>B�M��p.���׽[��Zc�cC����`7�{om��\)?���־{y�?LW�b�=��=Q|�>��?!D:?��d� 'J?�4?��??E�=�>�<��>�m1��� >
�>����f�վ�>��%�!�G� �=����������B�$'�����<I���`�>��>8ۨ>SWܽ<X��l�M?t��>�&��̎R�Ud>ۋ�=a��acz>	�>Z��=H6����>D��>�Ǫ?$��n(�Zv=̉>�ц��R�=��;tB?���f?�3?7x�<e¯>�YN�sg?ݴ/>�X=���=��N>�ѥ=�b�>��>l�?>�)>~��E�>���?��S?�쒾��> �;�x=�>�"!>��>t����'�>��v>k6��.����H�~n�1�΄�l�C���?N~�>w�Z>������>'y�>bBi>��������o�>I�4?����w&�>z�^�N>O�>ۏ?Z���uŨ���;?$��?6J��s=��{?Ѭ�>�?b=x�w�����aB��'�Jh�*C�ؘc?�J����<k��?�����X�;�Ҿ�q?*�?�Q?�����w_?N�D?�,:>���>Nd��xxf<�[^�?)u��֩>W����6���>�j�T?�T�?�V�����b8>��B=`ٿ��.�>�<?wK�_��=>LK?z�ۿ���<MS��v=l�e��1��v
P��;�>�����fA������c���� �+�1��0]��h����-?�ξ�-����b>=��>p6�>��������?�1�>#��ʳ���e�@ֆ�E�J�A;>��M�>
��_|K��i���-?է��Q�4�Zp�>� ?�߻>������Bш?0���\�=����7�>�xX?�Z�-��%R?+�><�>�}�jF���񾍬�>Ė	?O0 ?�<�jz4>�5@=7�ѿPJɼ���;�>�ω�i�%���:��-Y>�Z���F9�EJ����8�W?dQ���>�=?<���~<�=�C=�@�j�/�ne��$�2�\��>�糿�p������R�˙�>�~�8O�4>n>9�;�C��a">R�Y��砾�	o>=�J?�����;ڂQ?�'�>��*���!�|z><�F>����Ӥ��L�>&��>�/����
����E?-�a;��>aǊ>g�>q��?�u�7d?��?N�Ծ��?R9?�>�E�>e�*>'>d�'>PV���X�<I�;?OU5?ON>2�g���>�·>GBe�\��>�o��$܂?k�=��X���>�a���I��x��r�9?����p��=Ai?�����>屑<����W�������1����>C�@��כ���a��㷽f�Y�,"
<x������q�=�5S�)��>[�U�W>�о�'?p��>g�W>�7ľ����R?\����?��;��o����=O:?��,�q��5���Q>w��������E�u�?Pe>GL����8�<wՑ>���=���7$�O8=�u)=�J?���ͽ�k
?-B#�I��/������>�I�>:ek�Ꮎ�w�>�
 ����>f7�?Y�D<�C�?po�<8�8??��	UF?���>�G���
¾Ϋ��x>����L��<&e>��?H��=�����~���>��>�~c���]�Tv��M���d��>8�ҽ�H��V"?�"���=T�����>�78���
>��:����>���>��!�`���Ƈ>W��)�Y��6���x�>n'9��r���o�>=lz>�t������0>�W~?����������XA>��i>�J>M�?q^�cR>Nwb��m?K�Ҿ,2>�0a�:&�>/�'>��@��_r�D�D?1bž�=� >�>��J����$;=�q?Xt��"�=�BZ��w	?�?>��ľ�z$��Ñ���ھ�D�>�g� ܮ�~g=�m9?rK=;�i¯�"n>J�T>�J���ـ����>*��>;�?�Ҿ�R"?���7Uk�Lv�>��>E6�=r*��NO��}�>���>o���7���U?��6>���	M��쎷�������k���&��(߾�4��ܮN?��%��>��<B�>�H��o�%>&�/< ��>��5��>�9(�lOf�?v��[M�>5�=h����x�<�j>�@ۼ�R[��\�N��>|陾R�<>�\Y���*n�>����6>�ߣ��&=�>�u??z���G	 ���A?���>�r�@�>����E"���>~��5����?��=ۍ>)N�����>���E�	>��(�Jݷ>Ɍ>	��*�J�k>��>�� ?|��=O�l?�?�8�c���<�e�=�!���)�#`�=�J/��7	?���ƾ:=?���>ﴝ�尾��|�>NDs>��>�F�� ���y�=�=�R8�����>�>��V��>�T�>����>����/�y��>��C����9B�>����I�=1.��:
u��↾ڴp=?���.�>��=|І��:����_���?�o>��l�=\u�>�		?��q�]9;��N:\�>�X��G^7�����t�'�)�=�L�>0#�>p� �0Q'��{��*��P�1?�-����>�Ƴ=�Ge�;qD>�y�>�!?�h��n�>�� ��
a?PZ��/?8`D>WY�=fҾ���=*�>��>R��� �đ��_پ]�>�p���>'}���a?z�2��߳�! ���>[nc<t���%��?�?��ξgg�;���>�޾א�P�+��5?= ������Ҽ=�~>GE"�8G\=��5�H��> �b��8��u>/��=�#�� �3'���>ɵ���Ȼ�+��R�_? ���j|�Ƙ?8i�;�]�~Z�>��A���_Zp>�^1>=�)>�����=[��=l�=�k9�����Ԋ�>gT�>��O=U��>�`��P`�����6�Ҿ�~
>�[�=P�t<)E�>�Qy�B��>�Do���>椾ӯ?��?-�q��\�=���=l�=�f	�6�F=�5?��=����񽾲�>u��>�%�`K>��f���>ʸ1>j��=�Q�=���sD�>���;>��>��?&�c=ڭ�>�5���?�z����?���>�i==(V>�h&>�ǥ=�v>]Z&<Y'�=*`�>#֤�'򗽷�l=~�=$i]?DC�괚�PE�����`��Pu>O?���=�Z�Γ���?����XH�MT�@k?F#
><��\a�>��F��b+>n��>	�\�h���߳�R��>�-�=������>���=?y0>hNZ�ԑ�<Qo�=�MD��H�=��p=c�>4>���>_R3��C?$�=ɕL?C��XG?h��=��?&�����>��.=��_�������b�M�?�u=!�����D>������>�$#��g�>��S�]PW=�cq�	c ���%?�E�>c ��9�=���>M�>D��>x%h��#A��g���b?w�a����(>Q�R>˩��
=�Q�>2�>�Ծ��
�����5���>Ub�0�c>"OF���?B�}�}ߜ��?��	q"��F�>�Z<�������zw�`��&������=A�g=�(�>��3��X�>v\�A��<���������!?:A�>����c#=��=�U �@]�?�S��~`������T���#?D���M
>9Ez�pk�=��l��O���������>����8=��>%}�>�Ɍ>1���C���>��%=�i�S��+�?�
%='3=B�Ƚ�碾�v�)�����E��y>���>��:=��w�郲� e���vϽ�]>D��ۄ7�_z��4�Y�?5�>�b��ĸ	?�0�G=[ ���e?';����&>\��)�2?,�=.� >�W�:i�> �>.���y���>r�>��>tڷ���>V��<>8ﾂͅ>�ƨ=<"�͹�=Ǧ=�0���3>��&=�L>��N�m� �?�[���1����v�>���>�U��)����5��h�>���>q�p=�u�>���Jr�>�\>e��>�\��}?}�u>���TҽTT��sZ���/���5��ַ�{��<A��>Е^>E@̾��<$�>���=���Z[<��?� �>��5�
*>����Kć>=���5���>Z	K>�M�Ջ�>O1#�H�C�/�x=�=T!�>�;��Ǜ��U����>In>?�	�}�����8?I�ۺ��
>8�A� %�>�a��q��V&��n3?��t���>3r��� �>��>�[`<.HA�@?h�h>$6�>�r�����=��=�_��"�v�+��Ʒr>C�?Q?~�@?���=��F?�P>e`U?�ľ�'��@���!y��0�>��i>o���������Y?���v=޷
>�c�<6�9=��b���=
s�=lE>U�>�����>#
����Y>�g��&X=]��(��4�<����_�������>������U>{/�>GE�S�����>�9)?����P��j�f� �.>+5��1@��9 ?��-��=���>��~?�濾��ϽV��7?Q;���c����$���R����k1c>\��>I��<�X`�O����>Ic����t�/B���X?(�L=d5��bm�>���b͏>ͬ��?j�?�`��i%�cTʾC��>rWn�K����<�?�2��x;��9
�=eF�>vl�����>�%ӽ;﫾G@�;ǛJ> M�����Fm�>&_�=mQ'>'�?���	=(�>R��x��=�N����U�k��"�x��M���e>8���>8�>!Rþ V�>*���Ԏ=��/�-�پ�[?-��>�b�W���$*>Œ ?��?�-Ϛ>���:�P>e���'>/�B����>�4�����>���>��)P����@=�!�>�ͽp����Nh���?�?�+�O��I5?��(>lݽ�+���݅���<>� ?2�u�d���}�<P��=ғ��о\��>E)>K�J>�Ap�<�F�b�>��ξx>bA?��Y�>�U6��֝��w�=k�V>r<�M����>o̅>Ħ>Oý���W��>���kp�{�R�@�q�%�ʾ�9�='��=�b��-Խ�ޚ�!Hb?��ʾ:<�������.=���3͞�o��I�?��?����e�����<+�>9�V>�Vd��%����>.Lg=/�u������n�>r�U>�d�=��A��@2?sb�>��*>l�?$�-=fGԽ�	�>��>Ww�<�>ϫ<������?�Og�4U"�Ug�=w��>�y9�qӆ=Z���>��j>��L>��=�50?D<>�ğ��v����?O����>�����:�>�TȾ�����ن>{�i=�&�J��*P?J�Z}Ͼ鏘��lJ?�+þ�S�1�Z�,
��i��,��Y~�/m�>/�6����>�^2<}�;?�2[>�߼���|>W��=�{�?hP�>�5ݾ�0�ѫ�>R��=C�v>%ھ���>��/��2P?�F<�|�����>��-=��4cľ�th��j�>J�=�.��ފ>��뾐mE?(5<�f��)�>�+?~��ഽ�0�q�p?
`�i*c�����U?b>v?�k{��vd>�$?��-=�F�>�y=�ѝ�?P��>���-�??�?��=�g�=�>�e�>b�?;,�=�5�><��=u;�>�Q->��^> W�>'!�>`�D?�#�>�-��S�Tܾv*i�rG�>�y��V?Z�M�i�U?
y"=I�پg�4?���>�	N�����U�����>ݪŽ���`A���=# %�?[P?���>�ֽi���lі>*]�tآ���6�-�^>��?��	�JT��g$y�L�|��O?Q^g�9`�>�<D8��s?�G>��S�`T9?���>����p��F(���>o;�=�W>�?@D���_Z>j<7����>ݗn�%��>M��>'���+�=�&>�>!?B�?�B�����G�vC�����F~(�G1h�+{;�D>U�"=gW�ϧ@>��;?����x�=��5�e$]?�_�#(r�s@{�Fȼ�C�� ��!��;��W>�q%��!<� �<W�:�*Pžk}��)0?�:D�{퇽{��o)�>	��>�d������\��-ӾI�?T���Dn���v>^߽�_?�|v�`��8g5>��枹>���Pо�]�~P?���*���z>���>��k�U!	��z�?�S>)�0����"+h?�zr>�<�x��>�_?v�^��*�>���9�>CHG?���i�E?����C1�������n�?�<��f4�>h	��ל>��B���_k?/BZ>���X�P���`0�>��3�J]=���y>Vm�>�{?��>1��>�s�=]��;�l��|�=?-5�𖣾;����S���C�ľ<O ��I]=�+l>�����~�;�U>=���������Q�_?�)�C������Q*<�g>�hb>�n>��#?�'N����ꪉ�PR�+CO>:�?�_L��[�>"I>*����(?��*�Ϸf?m5?&d@��o�����e��>�V���B�>����.���^M?����[��
�>1%���z�>�3���$��\��>�Pg��X@�*�ؾt�%��\>犿r�3��=v�	����,C��1ѽ�^�?5'��<��a�.>-�Ͼ���>�p�>�hX���d>}��>�{�>�~?M����\?�t>�~s���Hd>�E>�H?�^2��vϾ �� �=u��t��ʾ�q���*?�c�-L�z���Ŭ:�XFT=ā���<��Vy?J����@>}4�&Ă�?�=��>�����l=��[>��>,��=O$�������J�>�G��/ྩ��>���> �����>�@�=�1?��->�q��$p�=y�P?´S>�ˑ>A��;���P�ս�FY��ck>�Λ�Ƕ�����<;f��asо�uq����>��4��R��E
޾GE�=�y�=���>>U��>!T>�~T��^þ��㾣W�>`8�=��=�f�p�?R?(oj����>�e? �?�8?D�p���=���E>v�?��>%A��z�? ˢ>Z�1��ZȽ�~q?�:�==	?�׭�M,��U�8?��нd}u�� %>q9��]?�)�.�}�n�]B�;�x��H�?"a> �w��L�>&�W>�	>�??�c=U8���>���\^=?��>�gd����@?�D�yZ�>�Jk������(?eR�0v>n;>������Q���%�v��=�p$=�H��
��>�U�ikk�DKC��_*?�Zk=/JE>�j���!?N��>�T:�/xF>���M=Q>���ő7>��6w�=K2�>v�>[�j����K��)�>Q�潺䉾���>G >�\-=���>�/�<��:>&w?l���(��	>�/?��\?��8>�*=f���D��E2��$���;'P��2�cx�0�=�;�ǽ��¾�7���<?�$�>b�w;�ʽ\�>�9�>`�c��'?f��;�RսV�#��1�>:�B7�>ٝ�=u�!�$w��@��J������Q���_�>�{G?�+����)�l�5���:X%���<<T-��Lh����Z�=��d>K�P?��0?U�>nM>���(T���ݼ:U;���"���i����,>�J�ܗ|���?�Υ=C�>Z��+l�=w\�=5�	����>]�=޸�>VI�?Vn�>5��>��[=��-��8꾲�U>�P�>�M��Q���)���[��n�>���>�1����>i���@C�>�l�>��a���>F�r>�p��v����7��:u�?	�>w������)�5c�g\����t��6�͟L>�=�j��BW�������>?}>.=�&>�ʽ�j,���Z?Ņ>���=�[;?�<?��7�Q:/>�!'>ڋ/>���?c�
z>��_�����M��>͏!>�m�>�(����>�þ"�?\����E?���>�i���K��n��'?�\��&ݾ6N@�H���;v>��=ӚӾz5�$�<��?���>��ľ1�= β��@>��A�b����� ?#�>ñ�=Ǆ�>��?��m>��=��>9�'�0n?�h��&y>���;c`���?6���#d�*�q=���=�#�>�ka>��U�z>�=N�� ���.�?6?ZG)?؍�*(>!?�Cx>���,�J�@I@>տ�� ۽y�=�|����?7ع>���XMs�ր�>SP>��<���h���Fu\?]0�����=�e�>:'��-�:�'>�2)>�v����ž�Y>/��=��X��/>pL�>>/?"��د�>aKI��6�>�>�=�����#�������&��LԾ��>g�A�����*]?t�6?�v<?K�>��?��?���>�E	>:h?>a�=���>q�;g8���F�H���s��	?���<���u�����=�� �\ݩ>3��Ӆb�j0����+���?���>���s�U�{J���4�1�0=����{�?,)>y5��W�K�˂s>ȑ��^g��q�>k3�>�?NT�������&2���%>�4����G8?�1�J���Zg?G�<���?�b��Á�ͷ4?����>3�Q��i���h�Kj��Ս<���<�����*�?�]z�C�%��[�LZ4?��>B>ח�v��>�,�>���=5޾��>@�Ѿ~�,�n��� 4^=	�?�k����@�')�>%�`�ٳX>���
����H�>�js�D��NՋ�5z�=��ѽ���>��v����=���>��>!nP��)���)��ߘz?��5�`zǾ}?�=��h��H5پ��@)����־���>�I��U�&p�>��ҽ�\�?L?��p��=�k�>p]��8S�g�>�Fվ���q���X>�D���҉>=Ô��x?��>�k����=�>[� ?҈�2��p,?>��>���=���v��>�,>ւ�>�7�]h[?
�??I?�0�5�=`#���S���}s�9��ҩֽY��=<8E>";h�#>o]>w��>E�M�#`Q���ݾM�u?������+UM�#	5=Iߞ=%HQ�����%?���Y��|s�>�Q>K�E�P�޼���2h?�=J������F�>V
���P��ؑ?犆�΍>��μ4:���Ll?WT��c��.2��f���=��o�qC���h?���>7R<��~��Yռ�K	>����%w>9�����>�؛�P.�"wF=*&�>�)Q�g>O��>g��>i ?x+q>��	?7^&?D�>�`&���H?ui�>O�>eQ�>|�d��#���Q���=q�c���?��>J1�>��">K9>��@��༷B�=T�?Ǩѽ��$;&�&�M)�>�j �5�`�*��=p��'@:<l�]��":>��K��%�ܖ>�>?G���*��Ծ��?"�=��WJ�D/�?+��3Rt��I���K�>Ts��ztǾ�֜��9��k�>PO��m4��`?[\M?{�3?չ�=�S}��E?>��d5�>�~\?��?�5�=aH$��>~7=\��=�.�>� 9�@1i��X����r�?t��6O�;��=e���$�=Zh)�m""��������w�
��"(���=�"�����p��+c>Ǥ>��T>J>X,`>�x>ݤ�>�	ۺ�h�>��>���>g�>�Y�>�J1���>��>70�>],>�@-?�=D>��><mU����>C�g><�>�i>���=]�5>�E��pv>�>=����½GY=�>	�i���H�>kἭ�6>6���ȺY�h��_��q:оF��<r��>;���E�=K��=��$�o�N����g��"���C����>����ǽ�T�*��>�0>���>X��
/�>��>P�'>���=e�>��)��
��ûa�J>��̾����=�>��>|N�8�\>#��>~��>uG>�4��w�=KXƾJ@�=��ļ��>F�:�;��>Jg�=��S>�B�=��������u>e9����=%���y�� 
�҄�>�'ҽ�����F>��<iB_�����>��=^T?DO=aq�h!;�|Gb;��>�]�<GPȽ|���n�����#?���>�JI���|�Kz��ͨ!�k�&+�<�a������2j|��GI�[� �%R�=T�ֽ�(�=>/E���������~M\��0�=��S�z����޾<mؼV�����Ӿ,E�=�X��& �9���Yt>��½�_���|�X8Q>S�>[�r:�=���)�����=W~�;&���?>��>ħ��G�H�.�<>_�}>^�y���G���>����;��]轈V��Z�>��׾������վ�;�QY���[�C���S=o� ����>�ES��0�>.,:��T�>�I?	A�>��n>�>
>h>վ0&��8�˯���8����<�Lݾ�>]Tۼ.s<�ҽ�����G���È>n9����׽X1�F�P>*���uV�����8�.>7��=�O<?�ʥ�x�V?@�>:�D>S咽��=�v+��|����j��Ku���i�w7Q�������=v�g�$�4��YF�#\>�܀�\$b=�=��o�L�`��}����;s2?amb��1�>h�=��?Ϸ���s��o��8�=��ľ�̏�:*������ث��W��\k���W>ֲ`��z�=�U��Htv��"_�p!>��>l��b@>YO�>�O>Q̾�{?hW�>KB�>Ma����>ݺ6>q�3>�T�XF!>�P���ȍ�i:�o�=�p���l>p?H?������Ћ���t>�]D���A�E^M�}�?��0>��M���>H:�>��>g�?W�Ƚr-�<��>��=1晽�\�J�^�1	=��ټm�����g�h�\[>���ΪN>ror>���>�R�����>�5=>��>�Bj�G K=&n�w'>+����P�=��g������4s>W%���Cj����=Q���j*������5>�l��v��\�n�,�n>�im�PE?o*\><�?�Y>Ў!>���<�ʺ�7������=��.?�S����!���>�u�>�A=�-8?���h2�=zV��f�=��<>�>?��>T����$>���>}��>�>yr�=�(�>�DB>��>˞�<�WL>��/��F�-�����[>�4!?c�+��=�-O>9�?Ƴ��Q��>4��>��>�`ľ��$;�8�>����\�>y�=��>��>P���A��y�Ľ��>�>�Ϣ��W�=��7���;֐;{��>=��=thf>q�<�y?��>%��>�=>�؊?j�?ݪ�<ܒ�>�_+?��>kKa;)H<< (>�9�:���&�=�����2>#��|�=M�!���K���*>\GN�`����==s���(��r��J�>y�<�/�o�ľ�J��2v���}="?(�7&>�m�>��z>�	�j�v��,��H�e>�ାe5��ph��w�`���m�=�(�y:�>7�b�ӻ4?��d>,��>���X�>Ғ��3t�>L>��~��a;�>��W>�q�=�5��<��襾d�w>�I��Qކ�_ʆ��>����g6*����1�>��	?ڠ\>�⍾V�M��> ��>$�_��W���>�K>
;���뾞�mjk>�c>�C�=9o�P7�k�X����R�=�^��i�"=!�r��d=?�->�Z�=et����>��̾�l���ľ���>o��=`�=�F����=�S> ����!��d���x� `�ڽJ?�iT�1O;�g�E�Q%�>m*=[4��)�B)?��/>s>R��hR��X�>�����{����>�D��<S���<���)���2=�{�H�p�o"���W=�Z0���½���Tn>,�ؾ�D������w=2�7�^3�>&%��[a��j4q>#���C�����7]>(q��)Y��˚�d ?��l��>�*6�=;?�2����=�L��x�>�~��+��<nDξ��>��Z>�eC��R���#8>G���%>�*K���>\۳�K��>���>�3?�[*��J��4�?+��>5��ʗ�_2[�z�O>*#��,{��^�g�,B0='�Q>�h'=Ȼ�����O�Ǿ1T>s5������@���ͽ���<{��<��F�H܎�Lǋ>0jھ��>�Q��+t�>��>�hо�{=�2>��>W���m�>���b�+>!X=�Fq�Fd�=�!=��H�&�Ӿ	;�������&�4�۾�=S�j��>��о�C�����xz?��?M�C��=u�K>f���t4
�^x�O!\>������M��A?�>|�+�:�����X�>�ؿ� �{>����`%?����QuX���A�q�ƾ 4�j�=K��=X)�\��m@ ������c>��>8��=l�j>+��>L'�>ba�>���>�H>���>���>zȽ�����4z>ag�����yb�>���=慍���ֽ%�>tн�&�=K.���E>�Q��@->��H�
>�>(����>�ͭ�����m���?ӽ��f���~ >X�?A0Q?ٕ]>�\�>8fX?�J1����&����g>����DU=L�?�>�Z>�[�>�RJ�>p���� =�P�q�>K_9�w�>�Y�<��?>̫X���=aR-��kS>�0����k>���<k��?���>�*>��=���??;:?�<���>)r-?�'@>t�>�&�R*>�<�pw�?��=u�?kB��tz>��X=�k�>�;y� ?<�3>o��>ܑ�Rs
>�����?��\
���x=�'8�ě3��*%��tͽ�mA��\�����R����'�\�-���ڽ��ؽ ў��m>"*wG���,�q_|����;�ui�
L�>�`��9\ �o2�>��<�8�!ˈ>����ɽ¯���f�mѐ��H>vv����>E >�Eo?ñQ=h�9����>T��>��z���=s��_�>�u�����X�V����>n'?�h��r�����K?�U��U={�6����>��%�� ��߽��%>��Ⱦ]c������#����M���򕽆��8��a�=O㦾��<�ǽ(��(B�<��5�)0=	���·3>�Q�r����e��I���6��&q�P�Խ����Ն澆^	�I^~=��sg���%7��3�=���4���^?���k�t���U4?�M#�`ja��֚��z2?$Έ�45�=�����>��>.>�Qɾ�\�~��4�!��
%��Ah�v��<B1᾽�Ѿ�t'>߯�=Q�Ѿp�=Zi�>�?\#>J>�y0>*��=�cļU�޼�>��~>ތ��
��|>N`�''��ʪ=\��>��?���=�EP>��3>�&]>�ھh۾:c>������D���>�&��3��[K>��&�����Dӽ�"3�Z�%�ȴ=[����I��0�y�J�e���G㾄���c�@�Ƽ�X���C�<>8x �j���I,�8mK}>|���K&�v�þe�>�}���ԏ�H� >l�P�~r>���>�'(?��Y;>a��>04A��~/��3�eΊ>B+>+C����ʾ2�v><>2r��v�K<.���0 A���^>h���_��=���>�E�=/R'�w��� j*��$1?��->U���~l��Q��>ڈ���c?����n����Q����=D5�=U쭼E����nF>��?!�_��4*?5�	?�i���!�>���<��>��g���k��7�>�B>G$(�i�<�x�>��~�[�l>_B�>�Q�>�Dd�Ͳ��)Ͼ0�������'�)�2>�b/>u�%?����>>������l>��	=����^�RǊ>�g�����>>ͽ(`x>P�>f�$?G[��վ�<�>3���.���$R:>�� ?v/���z�Q�C��'�=jWT=a��>Lj�>���?�%��)�=lU>*���R�����=���=�<��)��<�����]����t>4�O������>d�l�]A�<Y�==O�˽��g�Z��>���>!��>/�.=�`ܾ�餾v��o���a7?�Ƚ�5-��W�/�>A4>��̾���Q��>�k��A���׾.%'?��>u�ѽ�)��1�>U���[���O���˝>�I�=ы�����#?��׾Ģ���6��z)?�|�>iy��N�=��>�����n��嶾�G�f%>K���<��Nb�>p���s{�&7>=��������J��1>FY�><t���Ș<��<4�w>���>�5�C�"�T�x>C�O�7���㯾�@?Τ_�,E����<��x��=r >�T�TzQ�Ln��fl�=a܊=ᠪ=f �>�C�>��(�G`
�_�y��琾��Ծh�=gډ���=��?�����,>詫�����I=7U����c�켑Ė>������ �S>}�.>�
��z�>�sS?Sf%��eS=�ۋ=�_)��$�=5<�ތ���WB����>�9 �����b��>���>��Y=���ֆv>W��=LPY>�0ڽU��=���<���[��ݨԽ�&�>*��>Y8>�ϐ>ya��$>����]7���]>|y � ���������>��6���i=U�>>X�0��������A����pϾk�.>���F%>�@�e����(>ʤ?B0�̂?��+?��><hA��u;��2>-r|�x!�M'�=���=nv�>ٴ�=1@S���2��F<?քܽ����/Л<L?*v��oaH���~>�A>��@�)5���"�������>�K�=��<#��F�>���>?*j��Y�e I=��<�B������C�>���#i=���>t�sW���=� �>9-G��׾#7j���>�dB>�C'>h��>Щ�>gӽ�c��;�y���ƾr��;���=>�O>^�����=�T�=�6���\���潆/�=�!�=�C	�M⏾78>��< �ؾ�g���Y�{bJ>A���\=[�>���>�(c=�R�����ȓ>�x!�����>�^H�I읾�}>ǰ9��'>>F��Z>x
C�rD������@l����>_C�>;��>�+�>��g������� ��Y�E+��5?<tf�<�뽕G����'>`��>�ٽ\l���>��)>9��ƾp>V�=�w=pց�o�?�	n?@nI?�F¾��0=�f�<�n>}�N�A�L=f�>#	=����[<h׾�;˾�D�>)y1���i=E�K?�[��ۀ�>��)=�4�;]g�a4>E�>�>ý�����r�>d��>O�g>>@���I���+�>�6�>b�8��+S�l�><|!����ё�<���[J�ZF>��<@]��=G�����z�?_�>�1�P�$=p��=
^>/����9=���>~|ӽ{�P>p��]{�q��>� >ݷn>:��N� �e�T�R���޽�Fܽk�>�o5��T6��'>����.o�=Y�5<R|�����>�)�=��ӽ�� @g?L�l>�R�<F^H�W�-��ƻ��3������Ɵ�;i�����ϻx��w>�C�=D*����E>�����1��a�=[FJ�����_N>g��>�}��z�>���>J�=�:��G�{�Uq*����>��.��(���S�;�}>�=��<���>T��>�>��7}�������ٞ>�ƽ�NԾ���韋>���>뱎�⑆�m��= ��>D��=Ϡؾ��=G��m�~��Ċ��_�>7��=ڽM�z-�=��u<���څ�옆=�
���=�t?e�+G�<_R��1�>l��>R䳾��x=[:z�e�>��]i>m5��9�=��*�j>-]?>����=x�>�d/��G����i�b�=��>�R-�_���?�U�\��X�/�qLL?,+��������G��X���>{bk>J���Fq�=��[��#<�M����>�@�=�J�=��>v�=�����2�pƾ[�^>���>z|�=K>�>%���>�=k�=��?Pln������,������5P>f��<-?����>�Jp=0"w��*E>q?�����=9�ʾ��;�<��:��;<��"p���cQ>z�a��X��]�(>&������A?*8�=3rp��%:��j;>s���=������?�>/پ K��4��'�	>J�=�QL>�'�=`�E�� ?�n��?%�e�8�W`Z?w�>U��|����r�q0���/��:��r;ƾh->PE���9�=bV����潫��>�"?�9�|�y>唅>P�>PC4��=�!�>D�=g�����=���=�=�����j*���)=�7�����>y;V�r{�>&��>g�r�L/Խ��!<��n��T���k>�ȫ���>��O��b�=�9�!n�>�Ь�	e8�P����(�=��>R(#>E�(>�� >�#m�&�>�)���)�=��0�W�����I>���ֽ�"��M��Q�=�x�>o�>Y>$�>@hz>�x!���Ѻ��7?Q|ֽ�)=�R�>��Ddӽ�>�:@>��M�>�)�=<%���D>���;��>�R�=e=�����=��=�&��p.�(�G?��`�dɾV��=;���ۋ��ʶ�,(��s*���2v>D��>\��>�v�r����ve>�r?p4���>��>m6?�(�������6��X>(k�<�"&�`IX>w�=����ۼ�b{>�k[�u,�>��>�N�>�A�<-0j������ˮ���)���J���y>���{-U�4�:�ik�`i?���>�J�|��<n�=rC�=eh����
>Q��>�
��Y��6�׽چ�=�[پ״�=�j��G�->֣��#�:���=��>4H=�Յ��9^=�u���q>�ۃ��9(=��t>���=�#*>��������x>�f��d��Q_���a�>�,t�>辉�>��{P���y��\�U�(>����r����>�bԽ�v���4��=Wl���_>_y�>hw7��3M���v<����3�r��>%����6>�S�=R=��=pu�=���"-ݽ�:�=OEs>!�&>����>l�>N��=���X�
���>��>&����>���>��!>���*"��z=��#���Z>���q0��UP>�D>irZ>�
���q	
>��q��ʻ�3⩽͒�>��k�J�=(�V>��2���=<��>cc�=~f>�]㾾��&��>���=P�/=�ѽ@P�>�]v�S1����n��<�">��ݑ�>�C�n,����=��$?]�!��%Ž�3�>�<�;�/>��1�>{>Xp<�eD>�Z'��)%��n���j�>��>�ƾ�eC���=�,���ʾu!��>IP>{ee�U>W%?�����7=�,?���k��>�RU>44���>�=�=�h׾�)�>��7>���_>:|�>��=���=;��f�L>'�=!u����?��?�'�}���mf���P	?�>����݀a�f�>2g���=_�5�d^> x�=�����+���S?�bG�x;�������
?�z���N�r=������ ��gQ�,aw� �?��>ͳ�����y>I=dL?��>nHȾ�F�>	�>�lk>r�˾�.�=�'>��=k��>}�����E���>���>��U��������>K-�=�h����Q���=H	�>PK��L�      PK                      archive/data/8FB  fIž8�Z��jݾ�0ʾD�>�Pƾ���'��\�S�����V�+�Ĺ�g滾����_����S���XV=������Be�|)S�ٶ���žo�(�,=?>7��Y����1���7�X���u��I`�H�������G�Ҿ�<о2�)�����؊�|�6�u����z���oѾu���@� Y�5��,�˾dH���)I�0�ھr�e�rA��� �>۾�1�`��t�Ҿr�������		�����3˾�毾��*��0�+F��¾�M�������Kར	�ВվQ��"��Q��������d��(��ζ�|���Ӿ0�3�����2�����(���������<���G������� �X4̾�½_遾����ڋ�N���v��
�Ѿ��Ǿ�i����B��m������ ���x���W����a�A?��)�����I����ھ7�� R׾��w�M����'r�PK�,n      PK                      archive/data/9FB  ��c=�آ�)�?��S���=&��=K�
��V?e־5Ӽ9<��'F���b�/����>�AE=���>���>��?�@�>�����?oě>Hx�>,��;JѼ'�>o"?ry>��Ἳ<���?�?�>^�о%~
�qH`��$4?�WǾhG?>z��>��U��c��+p����>�Ɲ>5��>n��>�81��}�>�)�>��?.��f��>L����5s>�f?/}
����>�U>�U<�>��>�n>��>�O&?��b>z�2>d��?%�=���>t2�<���,�v=L|m>��"=���>�(���<���>S{���w�>䊖�Oj^>k�<��=ˠ��Y!T?c�H>�Ջ>z�&�UF�>�EJ?J�>ל�Y-�0�>�&��+?~+�=~�> ��>)��>&U�>)ޚ>�G?J����Q��1M�yЇ?�QT>�/?�=z2��D��>3�?�e\>Ͻ�>��=�[�>=��>e�־�X�|�>㛽WK>�|>�Ld>����'?k��h�5=�T�>F��k�?᳠�_���E�>��>x<��4?�1Q>��?]�D��a�>�,S=�]�ɺξ�`�>I�	<���>�4���u��>���>�N7>ꈾB��I<ϽW��>
j�=�L
>�%#�>�eƾ�ђ� 0��%�>�����e�� 8�����ɘ�<�	�$����=���>v�>��>�fp�����y��'��>�����(?"��=��>��U>Q1�=��5�ӽ�>�}��E
�{D�>%A�>h*?�@���껳��=�<�G >3nw��$�,�	?��?���>D��;q�.?]s�=����ꏽ R?�W ��|�>n�=nܼ���X>�'�h*޽��?G{�`Rս��8��>b������>׊`��� �P߹����&?�>�+$�\=/�J(Ӿq)>մG����>t�����I�u>��?Z��>vŴ�+b>d��>���� r�>��Q>V���Ѐ?����,��>�c�����>@.�<�DK=o?�>Db�>��� >�1?�>M����='�>��
�(l�����@r�E��>�J���i�B��>w�d��屾�4�>��K�'�0=�¾�zY;���>� ?M����-T?~݄��z*>w_־��W��|�>�,?j`?�/?T��VAB�,�<>9r�[�Ծ�-�
>U�>1c�>B2=1���"?fW=��U�����ǯ>�!�>]�>3}?(�۾@׾R�Ǿ%�6>�շ���'�3���>��>ն�<���>�⑾�R�>ւ>G��>��^=Wn���'��=�>��'>�)�=��ͽ�?���0����Y>g�b>��$?Pɼ����P	?�#�><݅����>���>B!�°̼��+�Ea����>ml߾}�=|��P<??��V=z�<ҀK���k=�/?�BV^��>�>�@���0?�x?�%?��罵�v=��?qɾ+Ҿo ��� ;��{��٩�>B��>i��>W�BoG>��>�'�>Tr���Q�a��;n��>�ں>[�;>�|�>�2��6��>>ӽ	��>��м�=���>�9�>T>?4�
��	�>��V���.?K��>,�>8�>u�<�1�=hڽ����>�>�\>7���q�>{��疍�쎃���>�ɋ>���<>�����>�݆>?�1�J�3gI=1�>�ჽ��!�l�c��>O<�|?�r$?Jق>U����>��=�>&��>���u?�<'?���d��>��<��z>�Yz>*�(?}�1?ݝR>�0���������UI�>4Ir<[_��ψ���0�.��f��>=��>sֻ<:Z?B~6>�YP�%>,;?��
=�m>*�|�e>N�"��=Ƅ�>h)�>���>��������o�:>ڒ���F��վ%Y<>�=��>�G=d�Z?�B�>�f�>��>��ɾ�p��-Ç��G�����>g.?�">x�>`R��ߐ�Wyb>��0=��;<�eB���+>�k��6�{�B?)-y��͔>L>PK����      PK                     C archive/versionFB? ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ3
PKўgU      PK          ����                     archive/data.pklPK          IVRN �   �               R  archive/data/0PK          .��                   Д  archive/data/1PK          ��)o                   �  archive/data/10PK          �PX                   ��  archive/data/2PK          v�@�                   �  archive/data/3PK          
��                   P�  archive/data/4PK          ����                   ��  archive/data/5PK          Y��                   Л  archive/data/6PK          ��L�                   �  archive/data/7PK          �,n                   �� archive/data/8PK          ����                   О archive/data/9PK          ўgU                   � archive/versionPK,       -                             ��     PK    ��        PK        ��   